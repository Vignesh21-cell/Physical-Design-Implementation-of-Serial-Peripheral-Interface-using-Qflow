* NGSPICE file created from spi_top.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

.subckt spi_top vdd gnd wb_clk_i wb_rst_i wb_adr_i[0] wb_adr_i[1] wb_adr_i[2] wb_adr_i[3]
+ wb_adr_i[4] wb_dat_i[0] wb_dat_i[1] wb_dat_i[2] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5]
+ wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12]
+ wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[30] wb_dat_i[31] wb_sel_i[0] wb_sel_i[1]
+ wb_sel_i[2] wb_sel_i[3] wb_we_i wb_stb_i wb_cyc_i miso_pad_i wb_dat_o[0] wb_dat_o[1]
+ wb_dat_o[2] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8]
+ wb_dat_o[9] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15]
+ wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[30] wb_dat_o[31] wb_ack_o wb_err_o wb_int_o ss_pad_o[0] ss_pad_o[1] ss_pad_o[2]
+ ss_pad_o[3] ss_pad_o[4] ss_pad_o[5] ss_pad_o[6] ss_pad_o[7] ss_pad_o[8] ss_pad_o[9]
+ ss_pad_o[10] ss_pad_o[11] ss_pad_o[12] ss_pad_o[13] ss_pad_o[14] ss_pad_o[15] ss_pad_o[16]
+ ss_pad_o[17] ss_pad_o[18] ss_pad_o[19] ss_pad_o[20] ss_pad_o[21] ss_pad_o[22] ss_pad_o[23]
+ ss_pad_o[24] ss_pad_o[25] ss_pad_o[26] ss_pad_o[27] ss_pad_o[28] ss_pad_o[29] ss_pad_o[30]
+ ss_pad_o[31] sclk_pad_o mosi_pad_o
XFILL_9_6_0 gnd vdd FILL
XFILL_17_5_0 gnd vdd FILL
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_360 BUFX4_156/Y AOI21X1_90/B AOI21X1_90/Y gnd AOI22X1_41/C vdd OAI21X1
XOAI21X1_382 BUFX4_156/Y OAI21X1_382/B OAI21X1_382/C gnd AOI22X1_49/C vdd OAI21X1
XOAI21X1_371 INVX2_60/Y MUX2X1_29/S OAI21X1_613/C gnd OAI21X1_371/Y vdd OAI21X1
XOAI21X1_393 BUFX4_156/Y OAI21X1_393/B OAI21X1_393/C gnd AOI22X1_53/C vdd OAI21X1
XFILL_23_3_0 gnd vdd FILL
XMUX2X1_28 MUX2X1_38/A MUX2X1_28/B MUX2X1_28/S gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_39 wb_dat_i[3] INVX1_95/A MUX2X1_47/S gnd MUX2X1_39/Y vdd MUX2X1
XMUX2X1_17 wb_dat_i[30] MUX2X1_17/B BUFX4_90/Y gnd MUX2X1_17/Y vdd MUX2X1
XFILL_6_4_0 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XOAI21X1_190 INVX8_10/A OR2X2_1/A OR2X2_1/B gnd OAI21X1_191/C vdd OAI21X1
XDFFSR_9 INVX2_2/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XNAND2X1_21 BUFX4_19/Y wb_dat_i[12] gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_43 AOI21X1_9/Y NOR2X1_10/Y gnd DFFSR_73/D vdd NAND2X1
XNAND2X1_10 MUX2X1_29/S wb_dat_i[17] gnd OAI21X1_19/C vdd NAND2X1
XNAND2X1_32 BUFX4_111/Y wb_dat_i[7] gnd OAI21X1_91/C vdd NAND2X1
XNAND2X1_76 INVX8_9/A OR2X2_1/B gnd OAI22X1_49/B vdd NAND2X1
XNAND2X1_87 OR2X2_7/B NOR2X1_54/A gnd NOR2X1_49/B vdd NAND2X1
XNAND2X1_98 BUFX4_181/Y INVX1_91/Y gnd NAND2X1_98/Y vdd NAND2X1
XNAND2X1_65 MUX2X1_17/B BUFX4_113/Y gnd NAND3X1_86/A vdd NAND2X1
XNAND2X1_54 INVX1_94/A BUFX4_113/Y gnd NAND3X1_75/A vdd NAND2X1
XAOI22X1_41 MUX2X1_8/B BUFX4_250/Y AOI22X1_41/C AOI22X1_41/D gnd DFFSR_237/D vdd AOI22X1
XAOI21X1_214 INVX2_71/Y OAI21X1_686/B BUFX4_257/Y gnd OAI21X1_686/C vdd AOI21X1
XAOI22X1_30 BUFX4_98/Y INVX1_7/A INVX2_103/A BUFX4_69/Y gnd NAND3X1_86/B vdd AOI22X1
XAOI21X1_203 INVX8_23/A OAI21X1_580/Y BUFX4_7/Y gnd AOI22X1_81/D vdd AOI21X1
XAOI22X1_52 MUX2X1_8/A BUFX4_250/Y AOI22X1_52/C AOI22X1_52/D gnd DFFSR_221/D vdd AOI22X1
XAOI22X1_85 INVX2_75/Y BUFX4_145/Y AOI22X1_85/C AOI22X1_85/D gnd DFFSR_203/D vdd AOI22X1
XAOI22X1_63 INVX2_138/Y BUFX4_143/Y AOI22X1_63/C AOI22X1_63/D gnd DFFSR_200/D vdd
+ AOI22X1
XAOI22X1_74 INVX2_107/Y BUFX4_7/Y AOI22X1_74/C AOI22X1_74/D gnd DFFSR_162/D vdd AOI22X1
XNAND3X1_229 BUFX4_207/Y NAND3X1_229/B NAND3X1_229/C gnd AOI21X1_55/A vdd NAND3X1
XNAND3X1_207 MUX2X1_42/B BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_209/B vdd NAND3X1
XNAND3X1_218 INVX1_118/Y BUFX4_47/Y BUFX4_141/Y gnd NAND3X1_220/B vdd NAND3X1
XOAI22X1_3 INVX8_5/A INVX1_20/Y INVX8_2/A INVX2_23/Y gnd OAI22X1_3/Y vdd OAI22X1
XFILL_30_6_1 gnd vdd FILL
XDFFSR_205 INVX2_82/A DFFSR_70/CLK BUFX4_15/Y vdd DFFSR_205/D gnd vdd DFFSR
XDFFSR_216 INVX1_32/A CLKBUF1_52/Y BUFX4_16/Y vdd DFFSR_216/D gnd vdd DFFSR
XDFFSR_249 INVX4_7/A CLKBUF1_37/Y BUFX4_15/Y vdd DFFSR_249/D gnd vdd DFFSR
XDFFSR_227 INVX2_72/A CLKBUF1_15/Y BUFX4_18/Y vdd DFFSR_227/D gnd vdd DFFSR
XDFFSR_238 INVX2_115/A CLKBUF1_24/Y BUFX4_10/Y vdd DFFSR_238/D gnd vdd DFFSR
XFILL_21_6_1 gnd vdd FILL
XFILL_20_1_0 gnd vdd FILL
XINVX2_45 INVX2_45/A gnd INVX2_45/Y vdd INVX2
XINVX2_34 INVX2_34/A gnd INVX2_34/Y vdd INVX2
XINVX2_56 INVX2_56/A gnd MUX2X1_4/A vdd INVX2
XINVX2_23 OR2X2_8/B gnd INVX2_23/Y vdd INVX2
XINVX2_12 DFFSR_3/Q gnd INVX2_12/Y vdd INVX2
XINVX2_78 INVX2_78/A gnd INVX2_78/Y vdd INVX2
XINVX2_67 INVX2_67/A gnd INVX2_67/Y vdd INVX2
XFILL_29_7_1 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XINVX2_89 INVX2_89/A gnd INVX2_89/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XFILL_4_7_1 gnd vdd FILL
XOAI21X1_19 INVX1_10/Y BUFX4_187/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XNAND2X1_239 BUFX4_6/Y OAI21X1_644/Y gnd OAI21X1_646/C vdd NAND2X1
XNAND2X1_217 INVX4_12/A NOR2X1_195/Y gnd OAI21X1_558/B vdd NAND2X1
XNAND2X1_206 INVX8_17/A INVX1_146/Y gnd OAI21X1_446/B vdd NAND2X1
XNAND2X1_228 BUFX4_7/Y OAI21X1_613/Y gnd OAI21X1_616/C vdd NAND2X1
XBUFX4_190 wb_sel_i[2] gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_261 NOR2X1_261/A NOR2X1_261/B gnd NOR2X1_261/Y vdd NOR2X1
XNOR2X1_250 BUFX4_253/Y OR2X2_13/A gnd NOR2X1_250/Y vdd NOR2X1
XOAI21X1_701 BUFX4_124/Y INVX8_20/Y MUX2X1_48/Y gnd OAI21X1_702/C vdd OAI21X1
XBUFX4_85 BUFX4_85/A gnd MUX2X1_6/S vdd BUFX4
XBUFX4_63 BUFX4_66/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_41 BUFX4_45/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_52 INVX8_15/Y gnd BUFX4_52/Y vdd BUFX4
XBUFX4_96 INVX8_1/Y gnd BUFX4_96/Y vdd BUFX4
XBUFX4_30 INVX8_3/Y gnd BUFX4_30/Y vdd BUFX4
XBUFX4_74 BUFX4_76/A gnd BUFX4_74/Y vdd BUFX4
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_11 OR2X2_11/A OR2X2_13/B gnd OR2X2_11/Y vdd OR2X2
XXNOR2X1_6 OR2X2_4/Y INVX2_50/Y gnd OR2X2_6/A vdd XNOR2X1
XFILL_26_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX8_11 wb_rst_i gnd INVX8_11/Y vdd INVX8
XOAI21X1_553 MUX2X1_15/A BUFX4_24/Y OAI21X1_553/C gnd OAI21X1_554/B vdd OAI21X1
XINVX8_22 INVX8_22/A gnd INVX8_22/Y vdd INVX8
XOAI21X1_564 INVX2_143/Y BUFX4_20/Y OAI21X1_644/C gnd OAI21X1_565/B vdd OAI21X1
XOAI21X1_520 INVX2_116/Y BUFX4_87/Y OAI21X1_520/C gnd OAI21X1_520/Y vdd OAI21X1
XOAI21X1_542 NOR2X1_204/Y INVX2_93/Y BUFX4_151/Y gnd OAI21X1_542/Y vdd OAI21X1
XOAI21X1_531 INVX2_98/Y BUFX4_187/Y OAI21X1_605/C gnd OAI21X1_532/B vdd OAI21X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOAI21X1_575 INVX2_125/Y BUFX4_106/Y OAI21X1_575/C gnd OAI21X1_575/Y vdd OAI21X1
XOAI21X1_597 INVX4_10/A INVX8_22/Y INVX1_153/A gnd NOR2X1_235/B vdd OAI21X1
XOAI21X1_586 BUFX4_163/Y MUX2X1_19/Y OAI21X1_586/C gnd DFFSR_145/D vdd OAI21X1
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XOAI21X1_361 MUX2X1_8/B BUFX4_87/Y OAI21X1_522/C gnd AOI21X1_91/B vdd OAI21X1
XOAI21X1_383 MUX2X1_9/A BUFX4_20/Y OAI21X1_630/C gnd OAI21X1_383/Y vdd OAI21X1
XOAI21X1_394 INVX2_142/Y BUFX4_22/Y OAI21X1_644/C gnd OAI21X1_394/Y vdd OAI21X1
XOAI21X1_372 INVX2_121/Y BUFX4_188/Y OAI21X1_617/C gnd AND2X2_14/A vdd OAI21X1
XOAI21X1_350 BUFX4_155/Y AOI21X1_80/B AOI21X1_80/Y gnd AOI22X1_36/C vdd OAI21X1
XFILL_23_3_1 gnd vdd FILL
XMUX2X1_29 wb_dat_i[22] MUX2X1_29/B MUX2X1_29/S gnd MUX2X1_29/Y vdd MUX2X1
XMUX2X1_18 MUX2X1_42/A MUX2X1_18/B MUX2X1_18/S gnd MUX2X1_18/Y vdd MUX2X1
XFILL_6_4_1 gnd vdd FILL
XFILL_14_3_1 gnd vdd FILL
XOAI21X1_191 INVX8_10/A OR2X2_3/Y OAI21X1_191/C gnd DFFSR_99/D vdd OAI21X1
XOAI21X1_180 XNOR2X1_2/Y NOR2X1_46/B OAI21X1_180/C gnd DFFSR_109/D vdd OAI21X1
XAOI22X1_1 INVX8_6/Y NOR2X1_96/A NOR2X1_98/A INVX8_7/Y gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_77 AND2X2_4/Y AND2X2_5/Y gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_33 INVX1_17/A OAI22X1_47/C gnd OAI21X1_76/B vdd NAND2X1
XNAND2X1_44 NAND2X1_44/A NOR2X1_11/Y gnd DFFSR_74/D vdd NAND2X1
XNAND2X1_22 BUFX4_21/Y wb_dat_i[13] gnd OAI21X1_73/C vdd NAND2X1
XNAND2X1_55 INVX1_119/A BUFX4_116/Y gnd NAND3X1_76/A vdd NAND2X1
XNAND2X1_11 BUFX4_188/Y wb_dat_i[18] gnd OAI21X1_21/C vdd NAND2X1
XNAND2X1_66 INVX1_96/A BUFX4_113/Y gnd NAND3X1_87/A vdd NAND2X1
XFILL_28_1 gnd vdd FILL
XNAND2X1_88 INVX2_48/Y INVX1_88/A gnd OR2X2_4/A vdd NAND2X1
XNAND2X1_99 MUX2X1_3/Y BUFX4_63/Y gnd NAND2X1_99/Y vdd NAND2X1
XAOI22X1_20 BUFX4_99/Y INVX1_2/A INVX2_84/A BUFX4_68/Y gnd NAND3X1_81/B vdd AOI22X1
XAOI22X1_53 INVX2_142/Y BUFX4_247/Y AOI22X1_53/C AOI22X1_53/D gnd DFFSR_220/D vdd
+ AOI22X1
XAOI21X1_215 BUFX4_257/Y OAI21X1_687/Y BUFX4_4/Y gnd AOI22X1_86/D vdd AOI21X1
XAOI21X1_204 NOR2X1_244/Y BUFX4_153/Y OAI21X1_664/Y gnd OAI22X1_118/C vdd AOI21X1
XAOI22X1_75 INVX2_119/Y BUFX4_4/Y AOI22X1_75/C AOI22X1_75/D gnd DFFSR_158/D vdd AOI22X1
XAOI22X1_64 INVX2_123/Y BUFX4_143/Y AOI22X1_64/C AOI22X1_64/D gnd DFFSR_198/D vdd
+ AOI22X1
XAOI22X1_31 INVX8_6/Y INVX2_69/A INVX2_67/A INVX8_7/Y gnd NAND3X1_87/C vdd AOI22X1
XAOI22X1_42 INVX2_139/Y BUFX4_246/Y AOI22X1_42/C AOI22X1_42/D gnd DFFSR_236/D vdd
+ AOI22X1
XAOI22X1_86 INVX2_71/Y BUFX4_4/Y AOI22X1_86/C AOI22X1_86/D gnd DFFSR_163/D vdd AOI22X1
XNAND3X1_208 INVX2_126/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_209/C vdd NAND3X1
XNAND3X1_219 INVX2_135/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_220/C vdd NAND3X1
XOAI22X1_4 OAI22X1_4/A INVX1_22/Y INVX1_21/Y INVX8_7/A gnd NOR2X1_3/B vdd OAI22X1
XDFFSR_239 INVX2_57/A CLKBUF1_60/Y BUFX4_8/Y vdd DFFSR_239/D gnd vdd DFFSR
XDFFSR_217 INVX1_35/A CLKBUF1_45/Y BUFX4_17/Y vdd DFFSR_217/D gnd vdd DFFSR
XDFFSR_206 INVX2_117/A CLKBUF1_29/Y BUFX4_17/Y vdd DFFSR_206/D gnd vdd DFFSR
XDFFSR_228 INVX2_145/A CLKBUF1_10/Y BUFX4_9/Y vdd DFFSR_228/D gnd vdd DFFSR
XFILL_20_1_1 gnd vdd FILL
XINVX2_46 INVX2_46/A gnd INVX2_46/Y vdd INVX2
XINVX2_79 INVX2_79/A gnd MUX2X1_6/A vdd INVX2
XINVX2_35 INVX2_35/A gnd INVX2_35/Y vdd INVX2
XINVX2_57 INVX2_57/A gnd MUX2X1_4/B vdd INVX2
XINVX2_24 INVX4_3/A gnd INVX2_24/Y vdd INVX2
XINVX2_13 DFFSR_4/Q gnd INVX2_13/Y vdd INVX2
XINVX2_68 INVX2_68/A gnd INVX2_68/Y vdd INVX2
XFILL_28_2_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XNAND2X1_207 INVX8_17/A INVX1_147/Y gnd OAI21X1_458/B vdd NAND2X1
XNAND2X1_218 INVX4_12/A AND2X2_18/A gnd OAI21X1_566/B vdd NAND2X1
XNAND2X1_229 NOR2X1_224/Y MUX2X1_48/A gnd OAI21X1_615/C vdd NAND2X1
XBUFX4_180 INVX8_12/Y gnd BUFX4_180/Y vdd BUFX4
XBUFX4_191 NAND3X1_1/Y gnd OAI22X1_5/A vdd BUFX4
XNOR2X1_251 INVX8_25/Y NOR2X1_251/B gnd NOR2X1_251/Y vdd NOR2X1
XNOR2X1_240 INVX8_25/Y NOR2X1_240/B gnd MUX2X1_40/S vdd NOR2X1
XNOR2X1_262 NOR2X1_51/A INVX4_10/Y gnd NOR2X1_262/Y vdd NOR2X1
XOAI21X1_702 BUFX4_163/Y MUX2X1_47/Y OAI21X1_702/C gnd DFFSR_123/D vdd OAI21X1
XBUFX4_20 wb_sel_i[1] gnd BUFX4_20/Y vdd BUFX4
XBUFX4_86 wb_sel_i[3] gnd BUFX4_86/Y vdd BUFX4
XBUFX4_75 BUFX4_76/A gnd BUFX4_75/Y vdd BUFX4
XBUFX4_42 BUFX4_45/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_97 INVX8_1/Y gnd BUFX4_97/Y vdd BUFX4
XBUFX4_53 INVX8_15/Y gnd BUFX4_53/Y vdd BUFX4
XBUFX4_64 BUFX4_66/A gnd BUFX4_64/Y vdd BUFX4
XBUFX4_31 INVX8_3/Y gnd BUFX4_31/Y vdd BUFX4
XFILL_10_1 gnd vdd FILL
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XOR2X2_12 OR2X2_13/B OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XXNOR2X1_7 XOR2X1_5/A XOR2X1_5/B gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XINVX8_12 OR2X2_9/B gnd INVX8_12/Y vdd INVX8
XFILL_0_0_1 gnd vdd FILL
XINVX8_23 INVX8_23/A gnd INVX8_23/Y vdd INVX8
XOAI21X1_521 NOR2X1_197/Y MUX2X1_6/B BUFX4_148/Y gnd OAI21X1_521/Y vdd OAI21X1
XOAI21X1_598 MUX2X1_25/B NOR2X1_219/Y OAI21X1_598/C gnd MUX2X1_26/A vdd OAI21X1
XOAI21X1_554 BUFX4_149/Y OAI21X1_554/B MUX2X1_26/S gnd OAI22X1_113/D vdd OAI21X1
XOAI21X1_587 INVX4_10/A INVX8_22/Y INVX1_151/A gnd NOR2X1_232/B vdd OAI21X1
XOAI21X1_510 NOR2X1_190/Y INVX2_90/Y BUFX4_149/Y gnd OAI21X1_510/Y vdd OAI21X1
XOAI21X1_565 BUFX4_147/Y OAI21X1_565/B BUFX4_162/Y gnd OAI22X1_116/D vdd OAI21X1
XOAI21X1_576 NOR2X1_212/Y INVX2_95/Y BUFX4_147/Y gnd OAI21X1_576/Y vdd OAI21X1
XOAI21X1_543 INVX2_93/Y NAND2X1_9/B OAI21X1_621/C gnd OAI21X1_544/B vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XOAI21X1_532 BUFX4_151/Y OAI21X1_532/B BUFX4_161/Y gnd OAI22X1_109/D vdd OAI21X1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_384 BUFX4_156/Y OAI21X1_384/B OAI21X1_384/C gnd AOI22X1_50/C vdd OAI21X1
XOAI21X1_395 BUFX4_160/Y OAI21X1_395/B OAI21X1_395/C gnd AOI22X1_54/C vdd OAI21X1
XOAI21X1_340 INVX1_50/A NOR2X1_79/B BUFX4_171/Y gnd OAI22X1_81/A vdd OAI21X1
XOAI21X1_373 BUFX4_146/Y BUFX4_255/Y INVX2_121/A gnd OAI21X1_374/C vdd OAI21X1
XOAI21X1_351 INVX2_103/Y BUFX4_91/Y OAI21X1_508/C gnd AOI21X1_81/B vdd OAI21X1
XFILL_10_7_0 gnd vdd FILL
XOAI21X1_362 BUFX4_160/Y AOI21X1_92/B AOI21X1_92/Y gnd AOI22X1_42/C vdd OAI21X1
XMUX2X1_19 wb_dat_i[29] MUX2X1_19/B BUFX4_91/Y gnd MUX2X1_19/Y vdd MUX2X1
XAOI22X1_2 BUFX4_93/Y INVX1_9/A INVX2_145/A BUFX4_67/Y gnd AOI22X1_2/Y vdd AOI22X1
XOAI21X1_170 INVX8_10/Y OR2X2_1/A INVX2_44/A gnd OAI21X1_171/C vdd OAI21X1
XOAI21X1_181 AOI21X1_23/Y NOR2X1_44/Y NOR2X1_47/B gnd OAI21X1_182/C vdd OAI21X1
XOAI21X1_192 BUFX4_183/Y OR2X2_8/B INVX2_49/Y gnd OAI21X1_193/C vdd OAI21X1
XNAND2X1_78 AND2X2_5/A AND2X2_5/B gnd NOR3X1_1/C vdd NAND2X1
XNAND2X1_89 NAND2X1_89/A NOR2X1_49/B gnd NOR2X1_256/B vdd NAND2X1
XNAND2X1_67 wb_stb_i wb_cyc_i gnd NOR2X1_16/B vdd NAND2X1
XNAND2X1_45 NAND2X1_45/A NOR2X1_12/Y gnd DFFSR_75/D vdd NAND2X1
XNAND2X1_34 wb_adr_i[2] wb_adr_i[3] gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_12 BUFX4_190/Y wb_dat_i[19] gnd OAI21X1_23/C vdd NAND2X1
XNAND2X1_56 INVX1_105/A BUFX4_113/Y gnd NAND3X1_77/A vdd NAND2X1
XNAND2X1_23 BUFX4_23/Y wb_dat_i[14] gnd OAI21X1_45/C vdd NAND2X1
XAOI21X1_205 INVX2_72/Y OAI21X1_667/B BUFX4_267/Y gnd OAI21X1_667/C vdd AOI21X1
XAOI21X1_216 INVX2_74/Y OAI21X1_688/B BUFX4_260/Y gnd OAI21X1_688/C vdd AOI21X1
XAOI22X1_54 INVX2_112/Y BUFX4_247/Y AOI22X1_54/C AOI22X1_54/D gnd DFFSR_218/D vdd
+ AOI22X1
XAOI22X1_10 BUFX4_93/Y INVX1_13/A INVX2_136/A BUFX4_67/Y gnd NAND3X1_76/B vdd AOI22X1
XAOI22X1_65 INVX2_91/Y BUFX4_146/Y AOI22X1_65/C AOI22X1_65/D gnd DFFSR_197/D vdd AOI22X1
XAOI22X1_87 INVX2_74/Y BUFX4_3/Y AOI22X1_87/C AOI22X1_87/D gnd DFFSR_171/D vdd AOI22X1
XAOI22X1_32 BUFX4_98/Y INVX1_8/A INVX2_68/A BUFX4_70/Y gnd NAND3X1_87/B vdd AOI22X1
XAOI22X1_43 INVX2_109/Y BUFX4_248/Y AOI22X1_43/C AOI22X1_43/D gnd DFFSR_234/D vdd
+ AOI22X1
XAOI22X1_76 INVX2_113/Y BUFX4_7/Y AOI22X1_76/C AOI22X1_76/D gnd DFFSR_154/D vdd AOI22X1
XAOI22X1_21 INVX8_6/Y INVX2_116/A INVX2_117/A INVX8_7/Y gnd NAND3X1_82/C vdd AOI22X1
XFILL_24_6_0 gnd vdd FILL
XNAND3X1_209 BUFX4_64/Y NAND3X1_209/B NAND3X1_209/C gnd AOI21X1_51/B vdd NAND3X1
XOAI22X1_5 OAI22X1_5/A INVX2_11/Y INVX2_40/Y OAI22X1_5/D gnd NOR2X1_3/A vdd OAI22X1
XFILL_7_7_0 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XDFFSR_207 INVX2_59/A CLKBUF1_28/Y BUFX4_8/Y vdd DFFSR_207/D gnd vdd DFFSR
XDFFSR_218 INVX1_38/A CLKBUF1_41/Y BUFX4_17/Y vdd DFFSR_218/D gnd vdd DFFSR
XDFFSR_229 INVX2_92/A CLKBUF1_7/Y BUFX4_9/Y vdd DFFSR_229/D gnd vdd DFFSR
XINVX2_47 INVX2_47/A gnd INVX2_47/Y vdd INVX2
XINVX2_58 INVX2_58/A gnd MUX2X1_5/A vdd INVX2
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XINVX2_25 INVX4_4/A gnd INVX2_25/Y vdd INVX2
XINVX2_69 INVX2_69/A gnd INVX2_69/Y vdd INVX2
XINVX2_14 DFFSR_5/Q gnd INVX2_14/Y vdd INVX2
XFILL_30_4_0 gnd vdd FILL
XNAND2X1_219 INVX4_12/A AND2X2_19/A gnd OAI21X1_568/B vdd NAND2X1
XNAND2X1_208 INVX8_17/A INVX1_148/Y gnd OAI21X1_462/B vdd NAND2X1
XNOR2X1_263 INVX4_10/A INVX1_17/A gnd NOR2X1_263/Y vdd NOR2X1
XBUFX4_181 INVX8_12/Y gnd BUFX4_181/Y vdd BUFX4
XNOR2X1_241 INVX8_25/Y NOR2X1_241/B gnd MUX2X1_42/S vdd NOR2X1
XNOR2X1_252 INVX8_24/Y NOR2X1_253/B gnd NOR2X1_252/Y vdd NOR2X1
XNOR2X1_230 INVX8_25/Y NOR2X1_230/B gnd MUX2X1_32/S vdd NOR2X1
XBUFX4_170 NOR3X1_9/Y gnd INVX1_138/A vdd BUFX4
XBUFX4_192 NAND3X1_1/Y gnd OAI22X1_8/A vdd BUFX4
XOAI21X1_703 OR2X2_5/B INVX4_9/A BUFX4_123/Y gnd OAI22X1_121/D vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_4_5_0 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XBUFX4_43 BUFX4_45/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 wb_sel_i[1] gnd BUFX4_21/Y vdd BUFX4
XBUFX4_10 BUFX4_9/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_32 BUFX4_35/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_87 wb_sel_i[3] gnd BUFX4_87/Y vdd BUFX4
XBUFX4_76 BUFX4_76/A gnd BUFX4_76/Y vdd BUFX4
XBUFX4_98 INVX8_1/Y gnd BUFX4_98/Y vdd BUFX4
XBUFX4_54 INVX8_15/Y gnd BUFX4_54/Y vdd BUFX4
XBUFX4_65 BUFX4_66/A gnd BUFX4_65/Y vdd BUFX4
XFILL_10_2 gnd vdd FILL
XXNOR2X1_8 OR2X2_5/A INVX4_8/A gnd OR2X2_8/A vdd XNOR2X1
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XINVX8_13 INVX8_13/A gnd INVX8_13/Y vdd INVX8
XINVX8_24 INVX8_24/A gnd INVX8_24/Y vdd INVX8
XOAI21X1_555 NOR2X1_209/Y MUX2X1_2/A BUFX4_148/Y gnd OAI21X1_555/Y vdd OAI21X1
XOAI21X1_522 MUX2X1_6/B BUFX4_88/Y OAI21X1_522/C gnd OAI21X1_523/B vdd OAI21X1
XOAI21X1_588 INVX4_10/A INVX8_20/Y MUX2X1_22/Y gnd OAI21X1_589/C vdd OAI21X1
XOAI21X1_511 INVX2_90/Y BUFX4_91/Y OAI21X1_511/C gnd OAI21X1_512/B vdd OAI21X1
XOAI21X1_599 BUFX4_125/Y INVX8_22/Y INVX1_154/A gnd NOR2X1_236/B vdd OAI21X1
XOAI21X1_577 INVX2_95/Y MUX2X1_43/S OAI21X1_658/C gnd OAI21X1_578/B vdd OAI21X1
XOAI21X1_544 BUFX4_151/Y OAI21X1_544/B BUFX4_165/Y gnd OAI22X1_111/D vdd OAI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XOAI21X1_500 BUFX4_229/Y OAI21X1_500/B INVX8_16/A gnd OAI22X1_100/D vdd OAI21X1
XOAI21X1_533 BUFX4_126/Y INVX2_156/Y INVX1_146/Y gnd INVX1_155/A vdd OAI21X1
XOAI21X1_566 BUFX4_159/Y OAI21X1_566/B OAI21X1_566/C gnd AOI22X1_76/C vdd OAI21X1
XFILL_9_1 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XOAI21X1_341 BUFX4_178/Y MUX2X1_23/B BUFX4_34/Y gnd OAI22X1_82/A vdd OAI21X1
XOAI21X1_330 INVX2_106/A NOR2X1_89/B INVX1_138/A gnd OAI22X1_77/A vdd OAI21X1
XFILL_10_7_1 gnd vdd FILL
XAND2X2_8 OR2X2_5/A OR2X2_5/B gnd AND2X2_8/Y vdd AND2X2
XOAI21X1_385 MUX2X1_13/A BUFX4_22/Y OAI21X1_553/C gnd OAI21X1_385/Y vdd OAI21X1
XOAI21X1_352 BUFX4_156/Y AOI21X1_82/B AOI21X1_82/Y gnd AOI22X1_37/C vdd OAI21X1
XOAI21X1_396 INVX2_112/Y BUFX4_106/Y OAI21X1_567/C gnd OAI21X1_396/Y vdd OAI21X1
XOAI21X1_363 INVX2_139/Y BUFX4_89/Y OAI21X1_525/C gnd AOI21X1_93/B vdd OAI21X1
XOAI21X1_374 OAI21X1_374/A BUFX4_249/Y OAI21X1_374/C gnd DFFSR_230/D vdd OAI21X1
XFILL_9_4_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XOAI21X1_171 NOR2X1_46/B XNOR2X1_1/Y OAI21X1_171/C gnd DFFSR_105/D vdd OAI21X1
XOAI21X1_160 XOR2X1_1/A NOR2X1_46/B OAI21X1_160/C gnd DFFSR_100/D vdd OAI21X1
XOAI21X1_182 INVX1_73/Y NOR2X1_47/B OAI21X1_182/C gnd DFFSR_110/D vdd OAI21X1
XAOI22X1_3 INVX8_6/Y INVX2_93/A INVX2_91/A INVX8_7/Y gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_193 INVX1_83/Y BUFX4_183/Y OAI21X1_193/C gnd INVX1_107/A vdd OAI21X1
XNAND2X1_79 NOR2X1_43/B NOR2X1_25/Y gnd INVX8_10/A vdd NAND2X1
XNAND2X1_68 INVX1_75/A NOR2X1_22/Y gnd OR2X2_2/A vdd NAND2X1
XNAND2X1_46 NAND2X1_46/A NOR2X1_13/Y gnd DFFSR_76/D vdd NAND2X1
XNAND2X1_35 AOI21X1_1/Y NOR2X1_2/Y gnd DFFSR_65/D vdd NAND2X1
XNAND2X1_24 BUFX4_25/Y wb_dat_i[15] gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_57 MUX2X1_29/B BUFX4_116/Y gnd NAND3X1_78/A vdd NAND2X1
XNAND2X1_13 BUFX4_185/Y wb_dat_i[20] gnd OAI21X1_25/C vdd NAND2X1
XAOI21X1_206 BUFX4_267/Y OAI21X1_668/Y BUFX4_247/Y gnd AOI22X1_82/D vdd AOI21X1
XAOI21X1_217 BUFX4_258/Y OAI21X1_689/Y BUFX4_3/Y gnd AOI22X1_87/D vdd AOI21X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XAOI22X1_33 INVX1_67/Y NOR2X1_46/B NOR2X1_46/Y AOI22X1_33/D gnd DFFSR_112/D vdd AOI22X1
XAOI22X1_55 INVX2_100/Y BUFX4_247/Y AOI22X1_55/C AOI22X1_55/D gnd DFFSR_217/D vdd
+ AOI22X1
XAOI22X1_77 INVX2_101/Y BUFX4_4/Y AOI22X1_77/C AOI22X1_77/D gnd DFFSR_153/D vdd AOI22X1
XAOI22X1_66 INVX2_147/Y BUFX4_143/Y AOI22X1_66/C AOI22X1_66/D gnd DFFSR_196/D vdd
+ AOI22X1
XAOI22X1_11 INVX8_6/Y INVX2_98/A INVX2_99/A INVX8_7/Y gnd NAND3X1_77/C vdd AOI22X1
XAOI22X1_22 BUFX4_95/Y INVX1_3/A INVX2_115/A BUFX4_70/Y gnd NAND3X1_82/B vdd AOI22X1
XAOI22X1_88 INVX2_77/Y BUFX4_5/Y AOI22X1_88/C AOI22X1_88/D gnd DFFSR_155/D vdd AOI22X1
XAOI22X1_44 INVX2_97/Y BUFX4_245/Y AOI22X1_44/C AOI22X1_44/D gnd DFFSR_233/D vdd AOI22X1
XFILL_24_6_1 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 INVX8_5/A INVX1_23/Y INVX8_2/A INVX2_24/Y gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_7_7_1 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFSR_208 INVX2_130/A CLKBUF1_21/Y BUFX4_15/Y vdd DFFSR_208/D gnd vdd DFFSR
XDFFSR_219 INVX2_76/A CLKBUF1_40/Y BUFX4_17/Y vdd DFFSR_219/D gnd vdd DFFSR
XINVX2_26 INVX4_6/A gnd INVX2_26/Y vdd INVX2
XINVX2_15 DFFSR_6/Q gnd INVX2_15/Y vdd INVX2
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XINVX2_59 INVX2_59/A gnd MUX2X1_5/B vdd INVX2
XINVX2_37 INVX2_37/A gnd INVX2_37/Y vdd INVX2
XFILL_30_4_1 gnd vdd FILL
XNAND2X1_209 INVX8_19/A INVX1_145/Y gnd OAI21X1_465/B vdd NAND2X1
XBUFX4_182 INVX8_12/Y gnd NOR2X1_73/B vdd BUFX4
XNOR2X1_231 INVX8_25/Y NOR2X1_231/B gnd AND2X2_25/B vdd NOR2X1
XNOR2X1_220 INVX8_24/Y NOR2X1_236/B gnd MUX2X1_28/S vdd NOR2X1
XNOR2X1_242 INVX1_157/A BUFX4_154/Y gnd NOR2X1_242/Y vdd NOR2X1
XBUFX4_193 NAND3X1_1/Y gnd BUFX4_193/Y vdd BUFX4
XBUFX4_171 NOR3X1_9/Y gnd BUFX4_171/Y vdd BUFX4
XBUFX4_160 INVX8_14/Y gnd BUFX4_160/Y vdd BUFX4
XNOR2X1_253 INVX8_25/Y NOR2X1_253/B gnd MUX2X1_48/S vdd NOR2X1
XOAI21X1_704 INVX4_2/A INVX4_9/A BUFX4_123/Y gnd OAI22X1_122/D vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XFILL_29_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_4_5_1 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XFILL_12_4_1 gnd vdd FILL
XBUFX4_44 BUFX4_45/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_22 wb_sel_i[1] gnd BUFX4_22/Y vdd BUFX4
XBUFX4_33 BUFX4_35/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_66 BUFX4_66/A gnd BUFX4_66/Y vdd BUFX4
XBUFX4_77 NOR3X1_8/Y gnd BUFX4_77/Y vdd BUFX4
XBUFX4_55 INVX8_15/Y gnd BUFX4_55/Y vdd BUFX4
XBUFX4_11 BUFX4_9/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_88 wb_sel_i[3] gnd BUFX4_88/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_99 INVX8_1/Y gnd BUFX4_99/Y vdd BUFX4
XFILL_10_3 gnd vdd FILL
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XXNOR2X1_9 XNOR2X1_9/A INVX4_4/A gnd XNOR2X1_9/Y vdd XNOR2X1
XINVX2_160 NOR2X1_85/Y gnd INVX2_160/Y vdd INVX2
XOAI21X1_523 BUFX4_148/Y OAI21X1_523/B BUFX4_164/Y gnd OAI22X1_106/D vdd OAI21X1
XOAI21X1_512 BUFX4_147/Y OAI21X1_512/B BUFX4_162/Y gnd OAI22X1_103/D vdd OAI21X1
XOAI21X1_501 NOR2X1_184/Y INVX2_96/Y BUFX4_233/Y gnd OAI21X1_501/Y vdd OAI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XINVX8_14 INVX8_14/A gnd INVX8_14/Y vdd INVX8
XINVX8_25 INVX8_25/A gnd INVX8_25/Y vdd INVX8
XOAI21X1_556 MUX2X1_2/A BUFX4_25/Y OAI21X1_635/C gnd OAI21X1_557/B vdd OAI21X1
XOAI21X1_589 MUX2X1_26/S MUX2X1_21/Y OAI21X1_589/C gnd DFFSR_144/D vdd OAI21X1
XOAI21X1_578 BUFX4_150/Y OAI21X1_578/B BUFX4_166/Y gnd OAI22X1_117/D vdd OAI21X1
XOAI21X1_545 BUFX4_157/Y OAI21X1_545/B OAI21X1_545/C gnd AOI22X1_73/C vdd OAI21X1
XOAI21X1_534 BUFX4_157/Y OAI21X1_534/B OAI21X1_534/C gnd AOI22X1_71/C vdd OAI21X1
XOAI21X1_567 INVX2_113/Y MUX2X1_37/S OAI21X1_567/C gnd OAI21X1_567/Y vdd OAI21X1
XFILL_9_2 gnd vdd FILL
XNAND3X1_190 INVX2_117/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_191/C vdd NAND3X1
XFILL_26_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_320 NOR2X1_99/B INVX1_93/A BUFX4_33/Y gnd OAI22X1_74/A vdd OAI21X1
XOAI21X1_353 MUX2X1_9/B BUFX4_86/Y OAI21X1_511/C gnd AOI21X1_83/B vdd OAI21X1
XOAI21X1_342 NOR2X1_87/B INVX1_113/A BUFX4_37/Y gnd OAI22X1_82/D vdd OAI21X1
XOAI21X1_331 NOR2X1_78/B MUX2X1_17/B BUFX4_32/Y gnd OAI22X1_78/A vdd OAI21X1
XOAI21X1_364 BUFX4_155/Y AOI21X1_94/B AOI21X1_94/Y gnd AOI22X1_43/C vdd OAI21X1
XAND2X2_9 INVX1_88/Y AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XOAI21X1_386 BUFX4_156/Y OAI21X1_386/B OAI21X1_386/C gnd AOI22X1_51/C vdd OAI21X1
XOAI21X1_397 BUFX4_156/Y OAI21X1_397/B OAI21X1_397/C gnd AOI22X1_55/C vdd OAI21X1
XOAI21X1_375 BUFX4_158/Y OAI21X1_375/B OAI21X1_375/C gnd AOI22X1_47/C vdd OAI21X1
XFILL_9_4_1 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_172 NAND2X1_82/Y XNOR2X1_1/B NOR2X1_27/B gnd AND2X2_7/A vdd OAI21X1
XOAI21X1_161 INVX8_10/Y OR2X2_1/A INVX2_40/A gnd OAI21X1_162/C vdd OAI21X1
XOAI21X1_183 NOR3X1_2/Y AOI21X1_24/Y NOR2X1_47/B gnd NAND2X1_83/B vdd OAI21X1
XOAI21X1_194 INVX2_49/Y OR2X2_8/B XNOR2X1_3/Y gnd INVX1_85/A vdd OAI21X1
XAOI22X1_4 BUFX4_93/Y INVX1_10/A INVX2_92/A BUFX4_67/Y gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_150 BUFX4_28/Y BUFX4_120/Y INVX1_1/A gnd BUFX2_27/A vdd OAI21X1
XNAND2X1_25 wb_dat_i[0] MUX2X1_41/S gnd OAI21X1_77/C vdd NAND2X1
XNAND2X1_14 BUFX4_187/Y wb_dat_i[21] gnd OAI21X1_27/C vdd NAND2X1
XNAND2X1_69 INVX1_80/A NOR2X1_24/Y gnd OR2X2_2/B vdd NAND2X1
XNAND2X1_47 NAND2X1_47/A NOR2X1_14/Y gnd DFFSR_77/D vdd NAND2X1
XNAND2X1_36 AOI21X1_2/Y NOR2X1_3/Y gnd DFFSR_66/D vdd NAND2X1
XNAND2X1_58 INVX1_98/A BUFX4_116/Y gnd NAND3X1_79/A vdd NAND2X1
XAOI22X1_23 INVX8_6/Y INVX2_54/A INVX2_59/A INVX8_7/Y gnd NAND3X1_83/C vdd AOI22X1
XAOI21X1_207 INVX2_73/Y OAI21X1_669/B BUFX4_262/Y gnd OAI21X1_669/C vdd AOI21X1
XAOI22X1_12 BUFX4_98/Y INVX1_14/A INVX2_97/A BUFX4_69/Y gnd NAND3X1_77/B vdd AOI22X1
XAOI21X1_218 INVX2_77/Y OAI21X1_690/B INVX8_23/A gnd OAI21X1_690/C vdd AOI21X1
XAOI22X1_34 AOI22X1_34/A AOI22X1_34/B AOI22X1_34/C AOI22X1_34/D gnd BUFX4_228/A vdd
+ AOI22X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_3/C gnd NOR3X1_2/Y vdd NOR3X1
XAOI22X1_45 INVX2_136/Y BUFX4_244/Y AOI22X1_45/C AOI22X1_45/D gnd DFFSR_232/D vdd
+ AOI22X1
XAOI22X1_56 INVX2_133/Y BUFX4_248/Y AOI22X1_56/C AOI22X1_56/D gnd DFFSR_216/D vdd
+ AOI22X1
XAOI22X1_78 INVX2_134/Y BUFX4_7/Y AOI22X1_78/C AOI22X1_78/D gnd DFFSR_152/D vdd AOI22X1
XAOI22X1_67 INVX2_108/Y BUFX4_144/Y AOI22X1_67/C AOI22X1_67/D gnd DFFSR_194/D vdd
+ AOI22X1
XAOI22X1_89 INVX2_76/Y BUFX4_246/Y AOI22X1_89/C AOI22X1_89/D gnd DFFSR_219/D vdd AOI22X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_7/A INVX1_25/Y INVX1_24/Y OAI22X1_7/D gnd NOR2X1_4/B vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XDFFSR_209 INVX2_88/A CLKBUF1_60/Y BUFX4_8/Y vdd DFFSR_209/D gnd vdd DFFSR
XINVX2_49 OR2X2_5/A gnd INVX2_49/Y vdd INVX2
XINVX2_38 INVX2_38/A gnd INVX2_38/Y vdd INVX2
XINVX2_27 INVX2_52/A gnd INVX2_27/Y vdd INVX2
XINVX2_16 DFFSR_7/Q gnd INVX2_16/Y vdd INVX2
XCLKBUF1_1 CLKBUF1_7/A gnd CLKBUF1_1/Y vdd CLKBUF1
XBUFX4_150 INVX8_23/Y gnd BUFX4_150/Y vdd BUFX4
XBUFX4_161 INVX8_21/Y gnd BUFX4_161/Y vdd BUFX4
XBUFX4_172 BUFX4_179/A gnd NOR2X1_78/B vdd BUFX4
XOAI21X1_705 INVX4_7/A INVX4_9/A OAI21X1_705/C gnd OAI21X1_706/A vdd OAI21X1
XNOR2X1_254 OR2X2_8/B BUFX4_123/Y gnd NOR2X1_254/Y vdd NOR2X1
XNOR2X1_210 INVX4_12/Y INVX1_153/Y gnd NOR2X1_210/Y vdd NOR2X1
XNOR2X1_232 INVX8_25/Y NOR2X1_232/B gnd MUX2X1_34/S vdd NOR2X1
XBUFX4_183 INVX8_12/Y gnd BUFX4_183/Y vdd BUFX4
XBUFX4_194 NAND3X1_1/Y gnd INVX8_1/A vdd BUFX4
XNOR2X1_221 INVX8_24/Y NOR2X1_237/B gnd MUX2X1_30/S vdd NOR2X1
XNOR2X1_243 INVX8_25/Y NOR2X1_243/B gnd MUX2X1_44/S vdd NOR2X1
XFILL_28_0_1 gnd vdd FILL
XFILL_3_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XBUFX4_23 wb_sel_i[1] gnd BUFX4_23/Y vdd BUFX4
XBUFX4_89 wb_sel_i[3] gnd BUFX4_89/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_45 BUFX4_45/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_34 BUFX4_35/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_67 INVX8_5/Y gnd BUFX4_67/Y vdd BUFX4
XBUFX4_12 BUFX4_9/A gnd BUFX4_12/Y vdd BUFX4
XBUFX4_56 BUFX4_61/A gnd BUFX4_56/Y vdd BUFX4
XBUFX4_78 NOR3X1_8/Y gnd BUFX4_78/Y vdd BUFX4
XINVX2_150 INVX1_18/A gnd INVX2_150/Y vdd INVX2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XINVX8_26 wb_rst_i gnd BUFX4_9/A vdd INVX8
XOAI21X1_557 BUFX4_148/Y OAI21X1_557/B BUFX4_164/Y gnd OAI22X1_114/D vdd OAI21X1
XOAI21X1_513 NOR2X1_192/Y MUX2X1_15/B BUFX4_149/Y gnd OAI21X1_513/Y vdd OAI21X1
XFILL_22_7_0 gnd vdd FILL
XOAI21X1_524 NOR2X1_199/Y INVX2_140/Y BUFX4_147/Y gnd OAI21X1_524/Y vdd OAI21X1
XOAI21X1_502 INVX2_96/Y BUFX4_108/Y OAI21X1_658/C gnd OAI21X1_503/B vdd OAI21X1
XINVX8_15 INVX8_15/A gnd INVX8_15/Y vdd INVX8
XOAI21X1_535 INVX2_137/Y BUFX4_188/Y OAI21X1_609/C gnd OAI21X1_535/Y vdd OAI21X1
XOAI21X1_546 INVX2_146/Y BUFX4_185/Y OAI21X1_624/C gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_568 BUFX4_153/Y OAI21X1_568/B OAI21X1_568/C gnd AOI22X1_77/C vdd OAI21X1
XOAI21X1_579 BUFX4_159/Y OAI21X1_579/B OAI21X1_579/C gnd AOI22X1_81/C vdd OAI21X1
XFILL_13_7_0 gnd vdd FILL
XFILL_9_3 gnd vdd FILL
XNAND3X1_191 BUFX4_65/Y NAND3X1_191/B NAND3X1_191/C gnd AOI21X1_48/B vdd NAND3X1
XNAND3X1_180 INVX2_113/Y BUFX4_50/Y BUFX4_137/Y gnd NAND3X1_181/C vdd NAND3X1
XOAI21X1_354 BUFX4_156/Y AOI21X1_84/B AOI21X1_84/Y gnd AOI22X1_38/C vdd OAI21X1
XOAI21X1_321 NOR2X1_99/B INVX1_92/A BUFX4_38/Y gnd OAI22X1_74/D vdd OAI21X1
XOAI21X1_387 MUX2X1_4/A BUFX4_24/Y OAI21X1_635/C gnd OAI21X1_387/Y vdd OAI21X1
XOAI21X1_398 INVX2_100/Y BUFX4_108/Y OAI21X1_569/C gnd OAI21X1_398/Y vdd OAI21X1
XOAI21X1_343 OAI22X1_81/Y OAI22X1_82/Y INVX2_155/Y gnd OAI21X1_343/Y vdd OAI21X1
XOAI21X1_376 INVX2_92/Y BUFX4_190/Y OAI21X1_621/C gnd OAI21X1_376/Y vdd OAI21X1
XOAI21X1_365 INVX2_109/Y BUFX4_187/Y OAI21X1_528/C gnd AOI21X1_95/B vdd OAI21X1
XOAI21X1_332 BUFX4_178/Y MUX2X1_31/B BUFX4_36/Y gnd OAI22X1_78/D vdd OAI21X1
XOAI21X1_310 BUFX4_178/Y INVX1_96/A BUFX4_34/Y gnd OAI22X1_70/A vdd OAI21X1
XFILL_27_6_0 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XOAI21X1_173 INVX8_10/Y OR2X2_1/A INVX2_45/A gnd OAI21X1_174/C vdd OAI21X1
XOAI21X1_162 NOR2X1_46/B XOR2X1_1/Y OAI21X1_162/C gnd DFFSR_101/D vdd OAI21X1
XOAI21X1_184 INVX8_10/Y OR2X2_1/A INVX2_34/A gnd NAND2X1_83/A vdd OAI21X1
XOAI21X1_195 INVX1_85/Y NOR2X1_55/Y BUFX2_80/A gnd OAI21X1_196/C vdd OAI21X1
XOAI21X1_151 BUFX4_27/Y BUFX4_118/Y INVX1_2/A gnd BUFX2_28/A vdd OAI21X1
XAOI22X1_5 INVX8_6/Y INVX2_122/A INVX2_123/A INVX8_7/Y gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_140 BUFX4_31/Y BUFX4_120/Y INVX2_8/A gnd BUFX2_17/A vdd OAI21X1
XFILL_10_5_0 gnd vdd FILL
XNAND2X1_48 NAND2X1_48/A NOR2X1_15/Y gnd DFFSR_78/D vdd NAND2X1
XNAND2X1_26 MUX2X1_43/S wb_dat_i[1] gnd OAI21X1_79/C vdd NAND2X1
XNAND2X1_15 BUFX4_189/Y wb_dat_i[22] gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_37 AOI21X1_3/Y NOR2X1_4/Y gnd DFFSR_67/D vdd NAND2X1
XNAND2X1_59 MUX2X1_27/B BUFX4_114/Y gnd NAND3X1_80/A vdd NAND2X1
XNAND2X1_190 BUFX4_21/Y wb_dat_i[8] gnd OAI21X1_644/C vdd NAND2X1
XFILL_18_6_0 gnd vdd FILL
XAOI22X1_24 BUFX4_99/Y INVX1_4/A INVX2_57/A BUFX4_68/Y gnd NAND3X1_83/B vdd AOI22X1
XAOI22X1_13 INVX8_6/Y INVX2_110/A INVX2_111/A INVX8_7/Y gnd NAND3X1_78/C vdd AOI22X1
XAOI21X1_208 BUFX4_262/Y OAI21X1_670/Y BUFX4_248/Y gnd AOI22X1_83/D vdd AOI21X1
XAOI22X1_46 INVX2_60/Y BUFX4_244/Y AOI22X1_46/C AOI22X1_46/D gnd DFFSR_231/D vdd AOI22X1
XAOI22X1_57 INVX2_64/Y BUFX4_245/Y AOI22X1_57/C AOI22X1_57/D gnd DFFSR_215/D vdd AOI22X1
XAOI21X1_219 BUFX4_257/Y OAI21X1_691/Y BUFX4_5/Y gnd AOI22X1_88/D vdd AOI21X1
XAOI22X1_35 INVX2_68/Y BUFX4_246/Y AOI22X1_35/C AOI22X1_35/D gnd DFFSR_243/D vdd AOI22X1
XNOR3X1_3 NOR3X1_3/A OR2X2_2/A NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XAOI22X1_68 INVX2_135/Y BUFX4_144/Y AOI22X1_68/C AOI22X1_68/D gnd DFFSR_184/D vdd
+ AOI22X1
XAOI22X1_79 INVX2_65/Y BUFX4_3/Y AOI22X1_79/C AOI22X1_79/D gnd DFFSR_151/D vdd AOI22X1
XOAI22X1_8 OAI22X1_8/A INVX2_12/Y INVX2_41/Y OAI22X1_8/D gnd NOR2X1_4/A vdd OAI22X1
XAOI21X1_90 MUX2X1_8/B AOI21X1_90/B BUFX4_264/Y gnd AOI21X1_90/Y vdd AOI21X1
XFILL_19_1 gnd vdd FILL
XINVX2_28 NOR3X1_6/A gnd INVX2_28/Y vdd INVX2
XINVX2_39 INVX2_39/A gnd INVX2_39/Y vdd INVX2
XINVX2_17 DFFSR_8/Q gnd INVX2_17/Y vdd INVX2
XFILL_24_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A INVX4_9/A MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XFILL_15_4_0 gnd vdd FILL
XCLKBUF1_2 CLKBUF1_2/A gnd CLKBUF1_2/Y vdd CLKBUF1
XNOR2X1_233 INVX8_25/Y NOR2X1_233/B gnd AND2X2_26/B vdd NOR2X1
XBUFX4_162 INVX8_21/Y gnd BUFX4_162/Y vdd BUFX4
XNOR2X1_211 INVX4_12/Y INVX1_154/Y gnd NOR2X1_211/Y vdd NOR2X1
XBUFX4_173 BUFX4_179/A gnd NOR2X1_82/B vdd BUFX4
XBUFX4_184 wb_sel_i[2] gnd NAND2X1_9/B vdd BUFX4
XBUFX4_195 NOR2X1_1/Y gnd AND2X2_1/B vdd BUFX4
XNOR2X1_200 BUFX4_251/Y OR2X2_11/A gnd AND2X2_18/A vdd NOR2X1
XNOR2X1_222 INVX8_24/Y NOR2X1_238/B gnd AND2X2_22/B vdd NOR2X1
XBUFX4_151 INVX8_23/Y gnd BUFX4_151/Y vdd BUFX4
XBUFX4_140 BUFX4_142/A gnd BUFX4_140/Y vdd BUFX4
XOAI21X1_706 OAI21X1_706/A INVX4_10/Y OAI21X1_706/C gnd DFFSR_249/D vdd OAI21X1
XNOR2X1_255 INVX4_9/Y INVX1_84/Y gnd NOR2X1_255/Y vdd NOR2X1
XNOR2X1_244 OR2X2_13/B NOR2X1_247/B gnd NOR2X1_244/Y vdd NOR2X1
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XBUFX4_24 wb_sel_i[1] gnd BUFX4_24/Y vdd BUFX4
XBUFX4_68 INVX8_5/Y gnd BUFX4_68/Y vdd BUFX4
XBUFX4_57 BUFX4_61/A gnd BUFX4_57/Y vdd BUFX4
XBUFX4_13 BUFX4_9/A gnd BUFX4_13/Y vdd BUFX4
XBUFX4_35 BUFX4_35/A gnd BUFX4_35/Y vdd BUFX4
XBUFX4_46 OR2X2_6/Y gnd BUFX4_46/Y vdd BUFX4
XBUFX4_79 NOR3X1_8/Y gnd BUFX4_79/Y vdd BUFX4
XFILL_30_2_0 gnd vdd FILL
XINVX2_151 INVX2_151/A gnd INVX2_151/Y vdd INVX2
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XINVX2_140 INVX2_140/A gnd INVX2_140/Y vdd INVX2
XINVX8_16 INVX8_16/A gnd INVX8_16/Y vdd INVX8
XOAI21X1_514 MUX2X1_15/B BUFX4_92/Y OAI21X1_514/C gnd OAI21X1_515/B vdd OAI21X1
XFILL_22_7_1 gnd vdd FILL
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_503 BUFX4_234/Y OAI21X1_503/B BUFX4_41/Y gnd OAI22X1_101/D vdd OAI21X1
XOAI21X1_525 INVX2_140/Y BUFX4_89/Y OAI21X1_525/C gnd OAI21X1_526/B vdd OAI21X1
XOAI21X1_569 INVX2_101/Y BUFX4_111/Y OAI21X1_569/C gnd OAI21X1_569/Y vdd OAI21X1
XOAI21X1_558 BUFX4_153/Y OAI21X1_558/B OAI21X1_558/C gnd AOI22X1_75/C vdd OAI21X1
XOAI21X1_536 AND2X2_20/Y INVX2_61/Y BUFX4_151/Y gnd OAI21X1_536/Y vdd OAI21X1
XOAI21X1_547 BUFX4_159/Y OAI21X1_547/B OAI21X1_547/C gnd AOI22X1_74/C vdd OAI21X1
XFILL_29_3_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XOAI22X1_120 INVX2_78/Y BUFX4_45/Y OAI22X1_120/C OAI22X1_120/D gnd DFFSR_187/D vdd
+ OAI22X1
XNAND3X1_170 MUX2X1_32/B BUFX4_48/Y BUFX4_137/Y gnd NAND3X1_172/B vdd NAND3X1
XNAND3X1_192 INVX2_118/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_194/B vdd NAND3X1
XNAND3X1_181 BUFX4_205/Y NAND3X1_181/B NAND3X1_181/C gnd AOI21X1_47/A vdd NAND3X1
XOAI21X1_355 MUX2X1_13/B BUFX4_88/Y OAI21X1_514/C gnd AOI21X1_85/B vdd OAI21X1
XOAI21X1_322 OAI22X1_73/Y OAI22X1_74/Y INVX2_155/Y gnd OAI21X1_322/Y vdd OAI21X1
XOAI21X1_344 OAI21X1_344/A OAI21X1_344/B INVX2_157/A gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_388 INVX2_118/Y BUFX4_26/Y OAI21X1_638/C gnd AND2X2_16/A vdd OAI21X1
XOAI21X1_300 BUFX4_178/Y MUX2X1_27/B BUFX4_34/Y gnd OAI22X1_66/D vdd OAI21X1
XOAI21X1_311 BUFX4_178/Y INVX1_97/A BUFX4_36/Y gnd OAI22X1_70/D vdd OAI21X1
XOAI21X1_377 BUFX4_158/Y OAI21X1_377/B OAI21X1_377/C gnd AOI22X1_48/C vdd OAI21X1
XOAI21X1_399 BUFX4_155/Y OAI21X1_399/B OAI21X1_399/C gnd AOI22X1_56/C vdd OAI21X1
XOAI21X1_333 OAI22X1_77/Y OAI22X1_78/Y NOR2X1_72/Y gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_366 BUFX4_160/Y AOI21X1_96/B AOI21X1_96/Y gnd AOI22X1_44/C vdd OAI21X1
XDFFSR_190 INVX1_48/A CLKBUF1_35/Y BUFX4_17/Y vdd DFFSR_190/D gnd vdd DFFSR
XNAND3X1_1 wb_adr_i[4] wb_adr_i[3] INVX2_1/Y gnd NAND3X1_1/Y vdd NAND3X1
XFILL_27_6_1 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_2_6_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XOAI21X1_130 BUFX4_31/Y BUFX4_118/Y DFFSR_5/Q gnd BUFX2_7/A vdd OAI21X1
XOAI21X1_174 AND2X2_7/Y NOR2X1_46/B OAI21X1_174/C gnd DFFSR_106/D vdd OAI21X1
XOAI21X1_163 XOR2X1_1/A XOR2X1_1/B INVX1_68/A gnd AND2X2_6/B vdd OAI21X1
XOAI21X1_185 NAND2X1_84/Y NOR3X1_2/A NOR2X1_22/B gnd AOI22X1_33/D vdd OAI21X1
XOAI21X1_196 BUFX2_80/A INVX1_84/Y OAI21X1_196/C gnd INVX1_86/A vdd OAI21X1
XOAI21X1_152 BUFX4_28/Y BUFX4_120/Y INVX1_3/A gnd BUFX2_29/A vdd OAI21X1
XAOI22X1_6 BUFX4_93/Y INVX1_11/A INVX2_121/A BUFX4_67/Y gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_141 BUFX4_31/Y BUFX4_118/Y INVX2_9/A gnd BUFX2_18/A vdd OAI21X1
XNAND2X1_180 BUFX4_19/Y wb_dat_i[13] gnd OAI21X1_630/C vdd NAND2X1
XNAND2X1_38 AOI21X1_4/Y NOR2X1_5/Y gnd DFFSR_68/D vdd NAND2X1
XNAND2X1_191 INVX1_139/A NOR2X1_153/Y gnd OAI21X1_395/B vdd NAND2X1
XNAND2X1_16 NAND2X1_9/B wb_dat_i[23] gnd OAI21X1_31/C vdd NAND2X1
XNAND2X1_27 MUX2X1_35/S wb_dat_i[2] gnd OAI21X1_81/C vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_49 NAND2X1_49/A NAND2X1_49/B gnd DFFSR_79/D vdd NAND2X1
XFILL_18_6_1 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_25 INVX8_6/Y INVX2_132/A INVX2_130/A INVX8_7/Y gnd NAND3X1_84/C vdd AOI22X1
XAOI21X1_209 INVX2_69/Y OAI21X1_671/B BUFX4_259/Y gnd OAI21X1_671/C vdd AOI21X1
XAOI22X1_14 BUFX4_94/Y INVX1_15/A INVX2_109/A BUFX4_69/Y gnd NAND3X1_78/B vdd AOI22X1
XAOI22X1_47 INVX2_92/Y BUFX4_249/Y AOI22X1_47/C AOI22X1_47/D gnd DFFSR_229/D vdd AOI22X1
XAOI22X1_69 INVX2_150/Y BUFX4_143/Y AOI22X1_69/C AOI22X1_69/D gnd DFFSR_180/D vdd
+ AOI22X1
XAOI22X1_36 INVX2_103/Y BUFX4_244/Y AOI22X1_36/C AOI22X1_36/D gnd DFFSR_242/D vdd
+ AOI22X1
XAOI22X1_58 INVX2_124/Y BUFX4_248/Y AOI22X1_58/C AOI22X1_58/D gnd DFFSR_214/D vdd
+ AOI22X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XOAI22X1_9 INVX8_5/A INVX1_26/Y INVX8_2/A INVX2_25/Y gnd OAI22X1_9/Y vdd OAI22X1
XAOI21X1_91 BUFX4_264/Y AOI21X1_91/B BUFX4_250/Y gnd AOI22X1_41/D vdd AOI21X1
XAOI21X1_80 INVX2_103/Y AOI21X1_80/B BUFX4_262/Y gnd AOI21X1_80/Y vdd AOI21X1
XINVX2_29 XOR2X1_3/B gnd INVX2_29/Y vdd INVX2
XINVX2_18 INVX4_8/A gnd INVX2_18/Y vdd INVX2
XFILL_24_4_1 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_6/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_15_4_1 gnd vdd FILL
XCLKBUF1_3 CLKBUF1_3/A gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_31_1 gnd vdd FILL
XNOR2X1_256 INVX4_9/Y NOR2X1_256/B gnd NOR2X1_256/Y vdd NOR2X1
XBUFX4_152 INVX8_14/Y gnd BUFX4_152/Y vdd BUFX4
XBUFX4_174 BUFX4_179/A gnd NOR2X1_99/B vdd BUFX4
XBUFX4_196 NOR2X1_1/Y gnd AND2X2_2/B vdd BUFX4
XBUFX4_130 INVX8_4/Y gnd BUFX4_130/Y vdd BUFX4
XNOR2X1_212 INVX4_12/Y NOR2X1_226/B gnd NOR2X1_212/Y vdd NOR2X1
XBUFX4_163 INVX8_21/Y gnd BUFX4_163/Y vdd BUFX4
XNOR2X1_201 BUFX4_253/Y NOR2X1_201/B gnd AND2X2_19/A vdd NOR2X1
XNOR2X1_234 INVX8_25/Y NOR2X1_234/B gnd AND2X2_27/B vdd NOR2X1
XBUFX4_185 wb_sel_i[2] gnd BUFX4_185/Y vdd BUFX4
XNOR2X1_223 INVX8_24/Y NOR2X1_239/B gnd AND2X2_23/B vdd NOR2X1
XBUFX4_141 BUFX4_142/A gnd BUFX4_141/Y vdd BUFX4
XNOR2X1_245 NOR2X1_75/A INVX2_160/Y gnd NOR2X1_245/Y vdd NOR2X1
XOAI21X1_707 INVX2_48/A INVX4_9/A OAI21X1_707/C gnd OAI21X1_708/A vdd OAI21X1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XBUFX4_14 BUFX4_9/A gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 wb_sel_i[1] gnd BUFX4_25/Y vdd BUFX4
XBUFX4_58 BUFX4_61/A gnd BUFX4_58/Y vdd BUFX4
XBUFX4_69 INVX8_5/Y gnd BUFX4_69/Y vdd BUFX4
XBUFX4_47 OR2X2_6/Y gnd BUFX4_47/Y vdd BUFX4
XBUFX4_36 BUFX4_39/A gnd BUFX4_36/Y vdd BUFX4
XFILL_30_2_1 gnd vdd FILL
XINVX2_130 INVX2_130/A gnd MUX2X1_14/B vdd INVX2
XINVX2_152 NOR2X1_72/Y gnd NOR2X1_75/B vdd INVX2
XINVX2_141 INVX2_141/A gnd INVX2_141/Y vdd INVX2
XINVX8_17 INVX8_17/A gnd OR2X2_13/B vdd INVX8
XOAI21X1_515 BUFX4_149/Y OAI21X1_515/B MUX2X1_26/S gnd OAI22X1_104/D vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_526 BUFX4_150/Y OAI21X1_526/B BUFX4_166/Y gnd OAI22X1_107/D vdd OAI21X1
XOAI21X1_559 INVX2_119/Y BUFX4_26/Y OAI21X1_638/C gnd OAI21X1_559/Y vdd OAI21X1
XOAI21X1_537 INVX2_61/Y BUFX4_189/Y OAI21X1_613/C gnd OAI21X1_538/B vdd OAI21X1
XOAI21X1_504 BUFX4_158/Y OAI21X1_504/B OAI21X1_504/C gnd AOI22X1_69/C vdd OAI21X1
XOAI21X1_548 INVX2_107/Y BUFX4_22/Y OAI21X1_548/C gnd OAI21X1_548/Y vdd OAI21X1
XFILL_29_3_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XOAI22X1_121 INVX4_3/Y BUFX4_123/Y NOR2X1_255/Y OAI22X1_121/D gnd DFFSR_247/D vdd
+ OAI22X1
XOAI22X1_110 INVX2_61/Y BUFX4_161/Y OAI22X1_110/C OAI22X1_110/D gnd DFFSR_167/D vdd
+ OAI22X1
XNAND3X1_160 INVX1_107/A NAND3X1_160/B NAND3X1_160/C gnd NAND3X1_252/B vdd NAND3X1
XNAND3X1_193 INVX2_119/Y BUFX4_48/Y BUFX4_138/Y gnd NAND3X1_194/C vdd NAND3X1
XNAND3X1_182 MUX2X1_36/B BUFX4_47/Y BUFX4_136/Y gnd NAND3X1_184/B vdd NAND3X1
XNAND3X1_171 INVX2_108/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_172/C vdd NAND3X1
XOAI21X1_323 OAI21X1_323/A OAI21X1_323/B NOR2X1_74/Y gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_301 OAI22X1_65/Y OAI22X1_66/Y INVX2_155/Y gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_312 OAI22X1_69/Y OAI22X1_70/Y NOR2X1_72/Y gnd OAI21X1_312/Y vdd OAI21X1
XDFFSR_191 INVX2_58/A CLKBUF1_29/Y BUFX4_8/Y vdd DFFSR_191/D gnd vdd DFFSR
XOAI21X1_356 BUFX4_156/Y AOI21X1_86/B AOI21X1_86/Y gnd AOI22X1_39/C vdd OAI21X1
XOAI21X1_345 OAI21X1_345/A OAI21X1_345/B OR2X2_10/Y gnd BUFX4_277/A vdd OAI21X1
XDFFSR_180 INVX1_18/A CLKBUF1_7/A BUFX4_9/Y vdd DFFSR_180/D gnd vdd DFFSR
XOAI21X1_378 INVX2_145/Y BUFX4_185/Y OAI21X1_624/C gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_367 INVX2_97/Y BUFX4_189/Y OAI21X1_605/C gnd AOI21X1_97/B vdd OAI21X1
XOAI21X1_334 INVX2_109/A NOR2X1_71/A BUFX4_80/Y gnd OAI22X1_79/D vdd OAI21X1
XOAI21X1_389 BUFX4_144/Y BUFX4_253/Y INVX1_50/A gnd OAI21X1_390/C vdd OAI21X1
XNAND3X1_2 wb_we_i wb_stb_i wb_cyc_i gnd NOR2X1_1/B vdd NAND3X1
XFILL_26_1_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_164 INVX8_10/Y OR2X2_1/A INVX2_41/A gnd OAI21X1_165/C vdd OAI21X1
XOAI21X1_120 AND2X2_3/Y INVX2_44/Y NAND3X1_65/Y gnd DFFSR_52/D vdd OAI21X1
XOAI21X1_131 BUFX4_27/Y BUFX4_118/Y DFFSR_6/Q gnd BUFX2_8/A vdd OAI21X1
XOAI21X1_153 BUFX4_29/Y BUFX4_118/Y INVX1_4/A gnd BUFX2_30/A vdd OAI21X1
XOAI21X1_142 BUFX4_30/Y BUFX4_124/Y INVX1_9/A gnd BUFX2_19/A vdd OAI21X1
XAOI22X1_7 INVX8_6/Y INVX2_61/A INVX2_62/A INVX8_7/Y gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_175 INVX8_10/Y OR2X2_1/A INVX2_46/A gnd OAI21X1_176/C vdd OAI21X1
XOAI21X1_197 OR2X2_5/A OR2X2_5/B INVX4_2/A gnd NAND2X1_89/A vdd OAI21X1
XOAI21X1_186 NOR3X1_3/Y AOI21X1_25/Y NOR2X1_47/B gnd NAND2X1_85/B vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_181 NOR2X1_148/Y INVX1_139/A gnd OAI21X1_384/B vdd NAND2X1
XNAND2X1_17 wb_dat_i[8] BUFX4_19/Y gnd OAI21X1_93/C vdd NAND2X1
XNAND2X1_28 BUFX4_111/Y wb_dat_i[3] gnd OAI21X1_83/C vdd NAND2X1
XNAND2X1_170 BUFX4_187/Y wb_dat_i[18] gnd OAI21X1_617/C vdd NAND2X1
XNAND2X1_39 AOI21X1_5/Y NOR2X1_6/Y gnd DFFSR_69/D vdd NAND2X1
XNAND2X1_192 wb_dat_i[6] MUX2X1_41/S gnd OAI21X1_567/C vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XNOR3X1_5 OR2X2_7/B INVX4_7/Y OR2X2_7/A gnd NOR3X1_5/Y vdd NOR3X1
XAOI22X1_26 BUFX4_99/Y INVX1_5/A INVX2_128/A BUFX4_68/Y gnd NAND3X1_84/B vdd AOI22X1
XAOI22X1_37 MUX2X1_9/B BUFX4_243/Y AOI22X1_37/C AOI22X1_37/D gnd DFFSR_241/D vdd AOI22X1
XAOI22X1_59 INVX2_94/Y BUFX4_247/Y AOI22X1_59/C AOI22X1_59/D gnd DFFSR_213/D vdd AOI22X1
XAOI22X1_15 INVX8_6/Y INVX2_74/A INVX2_75/A INVX8_7/Y gnd NAND3X1_79/C vdd AOI22X1
XAOI22X1_48 INVX2_145/Y BUFX4_249/Y AOI22X1_48/C AOI22X1_48/D gnd DFFSR_228/D vdd
+ AOI22X1
XBUFX2_80 BUFX2_80/A gnd BUFX2_80/Y vdd BUFX2
XAOI21X1_70 NOR2X1_76/A NOR2X1_76/B NOR2X1_73/B gnd AOI22X1_34/C vdd AOI21X1
XAOI21X1_81 BUFX4_262/Y AOI21X1_81/B BUFX4_248/Y gnd AOI22X1_36/D vdd AOI21X1
XAOI21X1_92 INVX2_139/Y AOI21X1_92/B BUFX4_268/Y gnd AOI21X1_92/Y vdd AOI21X1
XINVX2_19 wb_adr_i[3] gnd INVX2_19/Y vdd INVX2
XXOR2X1_2 INVX4_7/A INVX4_6/A gnd XOR2X1_2/Y vdd XOR2X1
XFILL_6_0_1 gnd vdd FILL
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B MUX2X1_8/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 CLKBUF1_4/A gnd DFFSR_5/CLK vdd CLKBUF1
XBUFX4_120 DFFSR_245/Q gnd BUFX4_120/Y vdd BUFX4
XFILL_31_2 gnd vdd FILL
XNOR2X1_257 INVX4_9/Y INVX1_91/A gnd NOR2X1_257/Y vdd NOR2X1
XNOR2X1_235 INVX8_25/Y NOR2X1_235/B gnd AND2X2_28/B vdd NOR2X1
XBUFX4_164 INVX8_21/Y gnd BUFX4_164/Y vdd BUFX4
XBUFX4_131 INVX8_4/Y gnd BUFX4_131/Y vdd BUFX4
XBUFX4_142 BUFX4_142/A gnd BUFX4_142/Y vdd BUFX4
XBUFX4_153 INVX8_14/Y gnd BUFX4_153/Y vdd BUFX4
XNOR2X1_246 BUFX4_253/Y NOR2X1_247/B gnd NOR2X1_246/Y vdd NOR2X1
XBUFX4_186 wb_sel_i[2] gnd MUX2X1_29/S vdd BUFX4
XBUFX4_197 NOR2X1_1/Y gnd NAND3X1_9/A vdd BUFX4
XNOR2X1_213 BUFX4_176/Y INVX1_144/Y gnd INVX8_24/A vdd NOR2X1
XBUFX4_175 BUFX4_179/A gnd NOR2X1_96/B vdd BUFX4
XNOR2X1_202 BUFX4_253/Y NOR2X1_202/B gnd AND2X2_20/A vdd NOR2X1
XNOR2X1_224 INVX8_24/Y NOR2X1_240/B gnd NOR2X1_224/Y vdd NOR2X1
XOAI21X1_708 OAI21X1_708/A INVX4_10/Y OAI21X1_708/C gnd DFFSR_250/D vdd OAI21X1
XFILL_25_7_0 gnd vdd FILL
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XFILL_0_7_0 gnd vdd FILL
XBUFX4_15 BUFX4_9/A gnd BUFX4_15/Y vdd BUFX4
XBUFX4_26 wb_sel_i[1] gnd BUFX4_26/Y vdd BUFX4
XBUFX4_37 BUFX4_39/A gnd BUFX4_37/Y vdd BUFX4
XBUFX4_48 OR2X2_6/Y gnd BUFX4_48/Y vdd BUFX4
XBUFX4_59 BUFX4_61/A gnd BUFX4_59/Y vdd BUFX4
XFILL_16_7_0 gnd vdd FILL
XINVX2_131 INVX1_55/A gnd MUX2X1_15/A vdd INVX2
XINVX2_142 INVX1_44/A gnd INVX2_142/Y vdd INVX2
XINVX2_153 NOR2X1_74/Y gnd NOR2X1_75/A vdd INVX2
XINVX2_120 INVX1_48/A gnd INVX2_120/Y vdd INVX2
XINVX8_18 INVX8_18/A gnd INVX8_18/Y vdd INVX8
XOAI21X1_505 INVX2_150/Y MUX2X1_35/S OAI21X1_580/C gnd OAI21X1_506/B vdd OAI21X1
XOAI21X1_516 NOR2X1_194/Y MUX2X1_2/B BUFX4_149/Y gnd OAI21X1_516/Y vdd OAI21X1
XOAI21X1_549 NOR2X1_207/Y INVX2_89/Y BUFX4_147/Y gnd OAI21X1_549/Y vdd OAI21X1
XOAI21X1_527 AND2X2_18/Y INVX2_110/Y BUFX4_150/Y gnd OAI21X1_527/Y vdd OAI21X1
XOAI21X1_538 BUFX4_151/Y OAI21X1_538/B BUFX4_161/Y gnd OAI22X1_110/D vdd OAI21X1
XAOI21X1_190 NOR2X1_211/Y BUFX4_154/Y OAI21X1_563/Y gnd OAI22X1_116/C vdd AOI21X1
XOAI22X1_122 INVX4_4/Y BUFX4_123/Y NOR2X1_256/Y OAI22X1_122/D gnd DFFSR_248/D vdd
+ OAI22X1
XOAI22X1_111 INVX2_93/Y BUFX4_165/Y OAI22X1_111/C OAI22X1_111/D gnd DFFSR_165/D vdd
+ OAI22X1
XOAI22X1_100 INVX2_126/Y INVX8_16/A OAI22X1_100/C OAI22X1_100/D gnd DFFSR_182/D vdd
+ OAI22X1
XNAND3X1_150 INVX2_100/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_152/B vdd NAND3X1
XNAND3X1_194 BUFX4_207/Y NAND3X1_194/B NAND3X1_194/C gnd AOI21X1_49/A vdd NAND3X1
XNAND3X1_161 INVX2_103/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_163/B vdd NAND3X1
XNAND3X1_183 INVX2_114/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_184/C vdd NAND3X1
XNAND3X1_172 BUFX4_65/Y NAND3X1_172/B NAND3X1_172/C gnd AOI21X1_45/B vdd NAND3X1
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_302 OAI21X1_302/A OAI21X1_302/B INVX2_159/A gnd OAI21X1_302/Y vdd OAI21X1
XOAI21X1_324 INVX2_121/A BUFX4_222/Y BUFX4_79/Y gnd OAI22X1_75/D vdd OAI21X1
XOAI21X1_313 INVX2_73/A NOR2X1_71/A BUFX4_80/Y gnd OAI22X1_71/D vdd OAI21X1
XOAI21X1_335 INVX1_38/A NOR2X1_79/B INVX1_138/A gnd OAI22X1_79/A vdd OAI21X1
XOAI21X1_346 BUFX4_153/Y AOI21X1_78/B AOI21X1_78/Y gnd AOI22X1_35/C vdd OAI21X1
XDFFSR_192 INVX1_54/A CLKBUF1_28/Y BUFX4_8/Y vdd DFFSR_192/D gnd vdd DFFSR
XOAI21X1_357 MUX2X1_4/B BUFX4_90/Y OAI21X1_590/C gnd AOI21X1_87/B vdd OAI21X1
XDFFSR_181 INVX2_96/A CLKBUF1_19/Y BUFX4_10/Y vdd DFFSR_181/D gnd vdd DFFSR
XOAI21X1_368 BUFX4_158/Y AOI21X1_98/B AOI21X1_98/Y gnd AOI22X1_45/C vdd OAI21X1
XDFFSR_170 INVX2_110/A CLKBUF1_1/Y BUFX4_12/Y vdd DFFSR_170/D gnd vdd DFFSR
XOAI21X1_379 INVX2_106/Y BUFX4_26/Y OAI21X1_548/C gnd AND2X2_15/A vdd OAI21X1
XFILL_5_6_0 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XNAND3X1_3 AND2X2_1/B OAI21X1_1/Y BUFX4_95/Y gnd OAI21X1_2/C vdd NAND3X1
XOAI21X1_176 NOR2X1_46/B AOI21X1_22/Y OAI21X1_176/C gnd DFFSR_107/D vdd OAI21X1
XOAI21X1_165 NOR2X1_46/B AND2X2_6/Y OAI21X1_165/C gnd DFFSR_102/D vdd OAI21X1
XOAI21X1_187 INVX8_10/Y OR2X2_1/A INVX2_36/A gnd NAND2X1_85/A vdd OAI21X1
XOAI21X1_198 OR2X2_5/B INVX4_3/Y INVX1_85/A gnd NOR2X1_56/B vdd OAI21X1
XOAI21X1_154 BUFX4_29/Y INVX8_9/A INVX1_5/A gnd BUFX2_31/A vdd OAI21X1
XOAI21X1_110 AND2X2_3/Y INVX2_39/Y NAND3X1_60/Y gnd DFFSR_47/D vdd OAI21X1
XOAI21X1_132 BUFX4_27/Y INVX8_9/A DFFSR_7/Q gnd BUFX2_9/A vdd OAI21X1
XOAI21X1_121 INVX2_45/Y BUFX4_111/Y OAI21X1_89/C gnd NAND3X1_66/B vdd OAI21X1
XOAI21X1_143 BUFX4_30/Y BUFX4_124/Y INVX1_10/A gnd BUFX2_20/A vdd OAI21X1
XAOI22X1_8 BUFX4_98/Y INVX1_12/A INVX2_60/A BUFX4_69/Y gnd AOI22X1_8/Y vdd AOI22X1
XNAND2X1_182 BUFX4_21/Y wb_dat_i[12] gnd OAI21X1_553/C vdd NAND2X1
XNAND2X1_18 BUFX4_21/Y wb_dat_i[9] gnd OAI21X1_95/C vdd NAND2X1
XNAND2X1_193 INVX1_139/A NOR2X1_154/Y gnd OAI21X1_397/B vdd NAND2X1
XNAND2X1_160 NOR2X1_152/Y NOR2X1_71/Y gnd AOI21X1_92/B vdd NAND2X1
XNAND2X1_171 NOR2X1_157/Y NOR2X1_71/Y gnd INVX1_137/A vdd NAND2X1
XNAND2X1_29 MUX2X1_41/S wb_dat_i[4] gnd OAI21X1_85/C vdd NAND2X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_7/A vdd NOR3X1
XAOI22X1_38 MUX2X1_13/B BUFX4_250/Y AOI22X1_38/C AOI22X1_38/D gnd DFFSR_240/D vdd
+ AOI22X1
XAOI22X1_49 MUX2X1_9/A BUFX4_250/Y AOI22X1_49/C AOI22X1_49/D gnd DFFSR_225/D vdd AOI22X1
XAOI22X1_27 INVX8_6/Y INVX2_90/A INVX2_88/A INVX8_7/Y gnd NAND3X1_85/C vdd AOI22X1
XAOI22X1_16 BUFX4_93/Y INVX1_16/A INVX2_73/A BUFX4_67/Y gnd NAND3X1_79/B vdd AOI22X1
XBUFX2_81 INVX2_22/A gnd BUFX2_81/Y vdd BUFX2
XBUFX2_70 OR2X2_8/B gnd BUFX2_70/Y vdd BUFX2
XFILL_27_4_0 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XAOI21X1_60 INVX4_8/A INVX2_50/Y BUFX4_272/Y gnd AOI22X1_34/B vdd AOI21X1
XAOI21X1_71 INVX4_8/Y INVX1_91/A AOI21X1_71/C gnd NOR3X1_9/A vdd AOI21X1
XAOI21X1_82 MUX2X1_9/B AOI21X1_82/B BUFX4_267/Y gnd AOI21X1_82/Y vdd AOI21X1
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_93 BUFX4_265/Y AOI21X1_93/B BUFX4_246/Y gnd AOI22X1_42/D vdd AOI21X1
XFILL_18_4_0 gnd vdd FILL
XOAI22X1_90 INVX2_62/Y INVX8_16/A OAI22X1_90/C OAI22X1_90/D gnd DFFSR_199/D vdd OAI22X1
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_9/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 CLKBUF1_5/A gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_154 INVX8_14/Y gnd BUFX4_154/Y vdd BUFX4
XBUFX4_132 BUFX4_135/A gnd INVX8_7/A vdd BUFX4
XBUFX4_121 DFFSR_245/Q gnd BUFX4_121/Y vdd BUFX4
XBUFX4_143 INVX8_16/Y gnd BUFX4_143/Y vdd BUFX4
XBUFX4_110 wb_sel_i[0] gnd MUX2X1_37/S vdd BUFX4
XFILL_31_3 gnd vdd FILL
XNOR2X1_258 INVX4_9/Y INVX1_81/Y gnd NOR2X1_259/B vdd NOR2X1
XNOR2X1_236 INVX8_25/Y NOR2X1_236/B gnd AND2X2_29/B vdd NOR2X1
XBUFX4_198 NOR2X1_1/Y gnd NAND3X1_7/A vdd BUFX4
XFILL_17_1 gnd vdd FILL
XNOR2X1_247 INVX8_19/Y NOR2X1_247/B gnd NOR2X1_247/Y vdd NOR2X1
XBUFX4_187 wb_sel_i[2] gnd BUFX4_187/Y vdd BUFX4
XBUFX4_165 INVX8_21/Y gnd BUFX4_165/Y vdd BUFX4
XNOR2X1_225 INVX8_24/Y NOR2X1_241/B gnd AND2X2_24/B vdd NOR2X1
XBUFX4_176 BUFX4_179/A gnd BUFX4_176/Y vdd BUFX4
XNOR2X1_203 BUFX4_251/Y OR2X2_12/B gnd NOR2X1_203/Y vdd NOR2X1
XNOR2X1_214 INVX8_24/Y NOR2X1_230/B gnd MUX2X1_18/S vdd NOR2X1
XOAI21X1_709 OR2X2_4/B INVX4_9/A BUFX4_123/Y gnd OAI22X1_123/D vdd OAI21X1
XFILL_25_7_1 gnd vdd FILL
XFILL_0_7_1 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 INVX8_7/A gnd INVX8_7/Y vdd INVX8
XBUFX4_38 BUFX4_39/A gnd BUFX4_38/Y vdd BUFX4
XBUFX4_49 OR2X2_6/Y gnd BUFX4_49/Y vdd BUFX4
XBUFX4_27 INVX8_3/Y gnd BUFX4_27/Y vdd BUFX4
XBUFX4_16 BUFX4_9/A gnd BUFX4_16/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XFILL_16_7_1 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XINVX2_132 INVX2_132/A gnd MUX2X1_15/B vdd INVX2
XINVX2_110 INVX2_110/A gnd INVX2_110/Y vdd INVX2
XINVX2_121 INVX2_121/A gnd INVX2_121/Y vdd INVX2
XINVX2_143 INVX1_43/A gnd INVX2_143/Y vdd INVX2
XINVX2_154 INVX2_154/A gnd INVX2_154/Y vdd INVX2
XOAI21X1_517 MUX2X1_2/B BUFX4_86/Y OAI21X1_590/C gnd OAI21X1_518/B vdd OAI21X1
XOAI21X1_528 INVX2_110/Y MUX2X1_29/S OAI21X1_528/C gnd OAI21X1_529/B vdd OAI21X1
XOAI21X1_539 BUFX4_157/Y OAI21X1_539/B OAI21X1_539/C gnd AOI22X1_72/C vdd OAI21X1
XOAI21X1_506 BUFX4_146/Y OAI21X1_506/B BUFX4_244/Y gnd AOI22X1_69/D vdd OAI21X1
XINVX8_19 INVX8_19/A gnd INVX8_19/Y vdd INVX8
XAOI21X1_180 INVX2_146/Y OAI21X1_545/B BUFX4_258/Y gnd OAI21X1_545/C vdd AOI21X1
XAOI21X1_191 INVX2_113/Y OAI21X1_566/B INVX8_23/A gnd OAI21X1_566/C vdd AOI21X1
XOAI22X1_101 INVX2_96/Y BUFX4_42/Y OAI22X1_101/C OAI22X1_101/D gnd DFFSR_181/D vdd
+ OAI22X1
XOAI22X1_123 INVX2_51/Y BUFX4_123/Y NOR2X1_257/Y OAI22X1_123/D gnd DFFSR_251/D vdd
+ OAI22X1
XOAI22X1_112 INVX2_89/Y BUFX4_162/Y OAI22X1_112/C OAI22X1_112/D gnd DFFSR_161/D vdd
+ OAI22X1
XFILL_30_0_0 gnd vdd FILL
XNAND3X1_151 INVX2_101/Y BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_152/C vdd NAND3X1
XNAND3X1_140 BUFX4_63/Y NAND3X1_140/B NAND3X1_140/C gnd NAND3X1_141/C vdd NAND3X1
XNAND3X1_162 INVX2_104/Y BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_163/C vdd NAND3X1
XNAND3X1_173 INVX2_109/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_175/B vdd NAND3X1
XNAND3X1_184 BUFX4_64/Y NAND3X1_184/B NAND3X1_184/C gnd AOI21X1_47/B vdd NAND3X1
XNAND3X1_195 INVX1_113/Y BUFX4_48/Y BUFX4_138/Y gnd NAND3X1_197/B vdd NAND3X1
XFILL_22_5_1 gnd vdd FILL
XOAI21X1_347 INVX8_22/A INVX8_20/A INVX4_10/Y gnd BUFX4_45/A vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_369 INVX2_136/Y NAND2X1_9/B OAI21X1_609/C gnd AOI21X1_99/B vdd OAI21X1
XOAI21X1_303 INVX2_60/A BUFX4_222/Y BUFX4_79/Y gnd OAI22X1_67/D vdd OAI21X1
XOAI21X1_336 BUFX4_176/Y MUX2X1_29/B BUFX4_32/Y gnd OAI22X1_80/A vdd OAI21X1
XOAI21X1_325 INVX1_26/A BUFX4_222/Y BUFX4_169/Y gnd OAI22X1_75/A vdd OAI21X1
XOAI21X1_314 INVX2_76/A NOR2X1_71/A INVX1_138/A gnd OAI22X1_71/A vdd OAI21X1
XOAI21X1_358 BUFX4_160/Y AOI21X1_88/B AOI21X1_88/Y gnd AOI22X1_40/C vdd OAI21X1
XDFFSR_160 INVX1_55/A DFFSR_70/CLK BUFX4_14/Y vdd DFFSR_160/D gnd vdd DFFSR
XDFFSR_193 INVX2_87/A CLKBUF1_21/Y BUFX4_8/Y vdd DFFSR_193/D gnd vdd DFFSR
XBUFX4_1 BUFX4_7/A gnd BUFX4_1/Y vdd BUFX4
XDFFSR_171 INVX2_74/A CLKBUF1_52/Y BUFX4_16/Y vdd DFFSR_171/D gnd vdd DFFSR
XDFFSR_182 INVX1_24/A CLKBUF1_16/Y BUFX4_16/Y vdd DFFSR_182/D gnd vdd DFFSR
XFILL_29_1_0 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XFILL_5_6_1 gnd vdd FILL
XINVX4_1 wb_adr_i[4] gnd INVX4_1/Y vdd INVX4
XFILL_13_5_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_4 NAND3X1_7/A OAI21X1_3/Y BUFX4_99/Y gnd OAI21X1_4/C vdd NAND3X1
XOAI21X1_177 NOR2X1_43/Y NOR3X1_1/Y NOR2X1_47/B gnd OAI21X1_178/C vdd OAI21X1
XOAI21X1_188 NAND2X1_86/Y NOR3X1_3/A NOR2X1_23/B gnd AOI21X1_27/A vdd OAI21X1
XOAI21X1_166 INVX8_10/Y OR2X2_1/A INVX2_42/A gnd OAI21X1_167/C vdd OAI21X1
XOAI21X1_199 INVX1_87/Y NOR2X1_56/Y OR2X2_6/B gnd OAI21X1_200/C vdd OAI21X1
XOAI21X1_122 AND2X2_3/Y INVX2_45/Y NAND3X1_66/Y gnd DFFSR_53/D vdd OAI21X1
XOAI21X1_100 AND2X2_3/Y INVX2_34/Y NAND3X1_55/Y gnd DFFSR_58/D vdd OAI21X1
XOAI21X1_111 INVX2_40/Y BUFX4_106/Y OAI21X1_79/C gnd NAND3X1_61/B vdd OAI21X1
XOAI21X1_155 BUFX4_31/Y BUFX4_118/Y INVX1_6/A gnd BUFX2_32/A vdd OAI21X1
XOAI21X1_133 BUFX4_31/Y BUFX4_118/Y DFFSR_8/Q gnd BUFX2_10/A vdd OAI21X1
XAOI22X1_9 INVX8_6/Y INVX2_137/A INVX2_138/A INVX8_7/Y gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_144 BUFX4_30/Y BUFX4_124/Y INVX1_11/A gnd BUFX2_21/A vdd OAI21X1
XNAND2X1_19 BUFX4_23/Y wb_dat_i[10] gnd OAI21X1_97/C vdd NAND2X1
XNAND2X1_150 NOR2X1_147/Y NOR2X1_71/Y gnd AOI21X1_82/B vdd NAND2X1
XNAND2X1_161 BUFX4_88/Y wb_dat_i[24] gnd OAI21X1_525/C vdd NAND2X1
XNAND2X1_183 NOR2X1_149/Y INVX1_139/A gnd OAI21X1_386/B vdd NAND2X1
XNAND2X1_194 MUX2X1_43/S wb_dat_i[5] gnd OAI21X1_569/C vdd NAND2X1
XNAND2X1_172 INVX1_137/Y INVX8_14/A gnd NAND2X1_172/Y vdd NAND2X1
XAOI22X1_39 MUX2X1_4/B BUFX4_243/Y AOI22X1_39/C AOI22X1_39/D gnd DFFSR_239/D vdd AOI22X1
XAOI22X1_28 BUFX4_99/Y INVX1_6/A INVX2_86/A BUFX4_68/Y gnd NAND3X1_85/B vdd AOI22X1
XAOI22X1_17 INVX8_6/Y INVX2_140/A INVX2_141/A INVX8_7/Y gnd NAND3X1_80/C vdd AOI22X1
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XBUFX2_71 INVX4_3/A gnd BUFX2_71/Y vdd BUFX2
XBUFX2_60 DFFSR_89/Q gnd wb_dat_o[24] vdd BUFX2
XBUFX2_82 INVX8_3/A gnd BUFX2_82/Y vdd BUFX2
XFILL_27_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_72 AOI21X1_72/A AOI21X1_72/B NOR3X1_7/C gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_61 AOI21X1_61/A AOI21X1_61/B INVX4_6/Y gnd NOR2X1_70/B vdd AOI21X1
XAOI21X1_83 BUFX4_263/Y AOI21X1_83/B BUFX4_243/Y gnd AOI22X1_37/D vdd AOI21X1
XAOI21X1_50 AOI21X1_50/A AOI21X1_50/B BUFX4_81/Y gnd AOI21X1_50/Y vdd AOI21X1
XOAI21X1_1 INVX1_1/Y BUFX4_87/Y OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XAOI21X1_94 INVX2_109/Y AOI21X1_94/B BUFX4_261/Y gnd AOI21X1_94/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XFILL_18_4_1 gnd vdd FILL
XOAI22X1_91 INVX2_87/Y BUFX4_41/Y OAI22X1_91/C OAI22X1_91/D gnd DFFSR_193/D vdd OAI22X1
XOAI22X1_80 OAI22X1_80/A OAI22X1_80/B OAI22X1_80/C OAI22X1_80/D gnd OAI22X1_80/Y vdd
+ OAI22X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B MUX2X1_8/S gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 CLKBUF1_6/A gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_122 DFFSR_245/Q gnd INVX8_9/A vdd BUFX4
XNOR2X1_215 INVX8_24/Y NOR2X1_231/B gnd MUX2X1_20/S vdd NOR2X1
XBUFX4_166 INVX8_21/Y gnd BUFX4_166/Y vdd BUFX4
XBUFX4_177 BUFX4_179/A gnd NOR2X1_87/B vdd BUFX4
XBUFX4_133 BUFX4_135/A gnd BUFX4_133/Y vdd BUFX4
XBUFX4_188 wb_sel_i[2] gnd BUFX4_188/Y vdd BUFX4
XBUFX4_144 INVX8_16/Y gnd BUFX4_144/Y vdd BUFX4
XBUFX4_111 wb_sel_i[0] gnd BUFX4_111/Y vdd BUFX4
XBUFX4_155 INVX8_14/Y gnd BUFX4_155/Y vdd BUFX4
XNOR2X1_204 INVX4_11/Y NOR2X1_226/B gnd NOR2X1_204/Y vdd NOR2X1
XBUFX4_100 AND2X2_1/Y gnd OAI21X1_2/A vdd BUFX4
XFILL_31_4 gnd vdd FILL
XNOR2X1_259 INVX4_10/Y NOR2X1_259/B gnd NOR2X1_259/Y vdd NOR2X1
XFILL_17_2 gnd vdd FILL
XNOR2X1_237 INVX8_25/Y NOR2X1_237/B gnd MUX2X1_36/S vdd NOR2X1
XNOR2X1_248 INVX8_19/Y OR2X2_13/A gnd NOR2X1_248/Y vdd NOR2X1
XNOR2X1_226 BUFX4_259/Y NOR2X1_226/B gnd NOR2X1_226/Y vdd NOR2X1
XBUFX4_199 NOR2X1_1/Y gnd BUFX4_199/Y vdd BUFX4
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 wb_rst_i gnd INVX8_8/Y vdd INVX8
XBUFX4_17 BUFX4_9/A gnd BUFX4_17/Y vdd BUFX4
XBUFX4_28 INVX8_3/Y gnd BUFX4_28/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XBUFX4_39 BUFX4_39/A gnd BUFX4_39/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XINVX2_100 INVX1_35/A gnd INVX2_100/Y vdd INVX2
XINVX2_155 INVX2_155/A gnd INVX2_155/Y vdd INVX2
XINVX2_144 INVX1_42/A gnd INVX2_144/Y vdd INVX2
XINVX2_111 INVX2_111/A gnd INVX2_111/Y vdd INVX2
XINVX2_122 INVX2_122/A gnd INVX2_122/Y vdd INVX2
XINVX2_133 INVX1_32/A gnd INVX2_133/Y vdd INVX2
XOAI21X1_518 BUFX4_149/Y OAI21X1_518/B BUFX4_164/Y gnd OAI22X1_105/D vdd OAI21X1
XOAI21X1_507 AND2X2_17/Y INVX2_104/Y BUFX4_150/Y gnd OAI21X1_507/Y vdd OAI21X1
XOAI21X1_529 BUFX4_150/Y OAI21X1_529/B BUFX4_165/Y gnd OAI22X1_108/D vdd OAI21X1
XAOI21X1_170 NOR2X1_197/Y BUFX4_152/Y OAI21X1_521/Y gnd OAI22X1_106/C vdd AOI21X1
XAOI21X1_181 BUFX4_258/Y OAI21X1_546/Y BUFX4_1/Y gnd AOI22X1_73/D vdd AOI21X1
XAOI21X1_192 BUFX4_259/Y OAI21X1_567/Y BUFX4_5/Y gnd AOI22X1_76/D vdd AOI21X1
XOAI22X1_113 MUX2X1_15/A MUX2X1_26/S OAI22X1_113/C OAI22X1_113/D gnd DFFSR_160/D vdd
+ OAI22X1
XOAI22X1_102 INVX2_104/Y BUFX4_165/Y OAI22X1_102/C OAI22X1_102/D gnd DFFSR_178/D vdd
+ OAI22X1
XFILL_30_0_1 gnd vdd FILL
XNAND3X1_152 BUFX4_207/Y NAND3X1_152/B NAND3X1_152/C gnd NAND3X1_156/B vdd NAND3X1
XNAND3X1_141 INVX8_13/A NAND3X1_141/B NAND3X1_141/C gnd NAND3X1_142/C vdd NAND3X1
XNAND3X1_196 INVX2_120/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_197/C vdd NAND3X1
XNAND3X1_185 INVX2_66/Y OAI21X1_224/Y OAI21X1_225/Y gnd NAND3X1_211/B vdd NAND3X1
XNAND3X1_174 INVX2_110/Y BUFX4_46/Y BUFX4_141/Y gnd NAND3X1_175/C vdd NAND3X1
XNAND3X1_130 BUFX4_62/Y NAND3X1_130/B NAND3X1_130/C gnd NAND3X1_134/B vdd NAND3X1
XNAND3X1_163 BUFX4_206/Y NAND3X1_163/B NAND3X1_163/C gnd AOI21X1_44/A vdd NAND3X1
XDFFSR_161 INVX2_89/A CLKBUF1_29/Y BUFX4_8/Y vdd DFFSR_161/D gnd vdd DFFSR
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_348 BUFX4_125/Y INVX2_156/Y BUFX4_42/Y gnd BUFX4_250/A vdd OAI21X1
XOAI21X1_326 NOR2X1_96/B INVX1_114/A BUFX4_35/Y gnd OAI22X1_76/A vdd OAI21X1
XDFFSR_150 INVX1_25/A CLKBUF1_6/A BUFX4_16/Y vdd DFFSR_150/D gnd vdd DFFSR
XOAI21X1_315 BUFX4_176/Y INVX1_98/A BUFX4_32/Y gnd OAI22X1_72/A vdd OAI21X1
XOAI21X1_304 INVX2_64/A BUFX4_222/Y BUFX4_169/Y gnd OAI22X1_67/A vdd OAI21X1
XOAI21X1_337 NOR2X1_78/B MUX2X1_35/B BUFX4_39/Y gnd OAI22X1_80/D vdd OAI21X1
XOAI21X1_359 INVX2_115/Y BUFX4_92/Y OAI21X1_520/C gnd AOI21X1_89/B vdd OAI21X1
XDFFSR_172 INVX2_140/A CLKBUF1_45/Y BUFX4_17/Y vdd DFFSR_172/D gnd vdd DFFSR
XDFFSR_183 INVX2_63/A CLKBUF1_9/Y BUFX4_17/Y vdd DFFSR_183/D gnd vdd DFFSR
XBUFX4_2 BUFX4_7/A gnd BUFX4_2/Y vdd BUFX4
XDFFSR_194 INVX1_61/A CLKBUF1_54/Y BUFX4_9/Y vdd DFFSR_194/D gnd vdd DFFSR
XFILL_29_1_1 gnd vdd FILL
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd OR2X2_7/B vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 AND2X2_1/B OAI21X1_5/Y BUFX4_98/Y gnd OAI21X1_6/C vdd NAND3X1
XOAI21X1_101 INVX2_35/Y BUFX4_21/Y OAI21X1_71/C gnd NAND3X1_56/B vdd OAI21X1
XOAI21X1_112 AND2X2_3/Y INVX2_40/Y NAND3X1_61/Y gnd DFFSR_48/D vdd OAI21X1
XOAI21X1_189 NAND2X1_86/Y INVX1_80/Y NOR2X1_47/B gnd OAI22X1_50/C vdd OAI21X1
XOAI21X1_178 INVX1_71/Y NOR2X1_47/B OAI21X1_178/C gnd DFFSR_108/D vdd OAI21X1
XOAI21X1_167 NOR2X1_46/B AOI21X1_20/Y OAI21X1_167/C gnd DFFSR_103/D vdd OAI21X1
XOAI21X1_123 INVX2_46/Y MUX2X1_47/S OAI21X1_91/C gnd NAND3X1_67/B vdd OAI21X1
XOAI21X1_145 BUFX4_28/Y BUFX4_120/Y INVX1_12/A gnd BUFX2_22/A vdd OAI21X1
XOAI21X1_156 BUFX4_28/Y BUFX4_120/Y INVX1_7/A gnd BUFX2_33/A vdd OAI21X1
XOAI21X1_134 BUFX4_31/Y BUFX4_118/Y INVX2_2/A gnd BUFX2_11/A vdd OAI21X1
XNAND2X1_184 BUFX4_23/Y wb_dat_i[11] gnd OAI21X1_635/C vdd NAND2X1
XNAND2X1_140 OAI21X1_286/Y OAI21X1_291/Y gnd OAI21X1_302/A vdd NAND2X1
XNAND2X1_151 BUFX4_92/Y wb_dat_i[29] gnd OAI21X1_511/C vdd NAND2X1
XNAND2X1_195 INVX1_139/A NOR2X1_155/Y gnd OAI21X1_399/B vdd NAND2X1
XNAND2X1_173 NOR2X1_159/Y NOR2X1_71/Y gnd OAI21X1_375/B vdd NAND2X1
XNAND2X1_162 NOR2X1_71/Y NOR2X1_153/Y gnd AOI21X1_94/B vdd NAND2X1
XAOI22X1_29 INVX8_6/Y INVX2_104/A INVX2_105/A INVX8_7/Y gnd NAND3X1_86/C vdd AOI22X1
XAOI22X1_18 BUFX4_95/Y INVX1_1/A INVX2_139/A BUFX4_70/Y gnd NAND3X1_80/B vdd AOI22X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_9/A NOR3X1_9/C gnd NOR3X1_8/Y vdd NOR3X1
XOAI21X1_690 BUFX4_159/Y OAI21X1_690/B OAI21X1_690/C gnd AOI22X1_88/C vdd OAI21X1
XBUFX2_72 INVX4_4/A gnd BUFX2_72/Y vdd BUFX2
XBUFX2_61 DFFSR_90/Q gnd wb_dat_o[25] vdd BUFX2
XBUFX2_50 DFFSR_79/Q gnd wb_dat_o[14] vdd BUFX2
XAOI21X1_62 NOR2X1_70/A AOI21X1_62/B NOR2X1_70/B gnd AOI21X1_72/A vdd AOI21X1
XAOI21X1_73 AOI21X1_73/A AOI21X1_73/B NOR2X1_73/B gnd NOR3X1_9/C vdd AOI21X1
XAOI21X1_84 MUX2X1_13/B AOI21X1_84/B BUFX4_264/Y gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_95 BUFX4_262/Y AOI21X1_95/B BUFX4_248/Y gnd AOI22X1_43/D vdd AOI21X1
XOAI21X1_2 OAI21X1_2/A INVX1_1/Y OAI21X1_2/C gnd DFFSR_25/D vdd OAI21X1
XAOI21X1_51 AOI21X1_51/A AOI21X1_51/B INVX8_13/Y gnd AOI21X1_51/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XAOI21X1_40 AOI21X1_40/A AOI21X1_40/B INVX8_13/Y gnd AOI21X1_40/Y vdd AOI21X1
XOAI22X1_70 OAI22X1_70/A OAI22X1_70/B OAI22X1_70/C OAI22X1_70/D gnd OAI22X1_70/Y vdd
+ OAI22X1
XOAI22X1_92 MUX2X1_14/A BUFX4_44/Y OAI22X1_92/C OAI22X1_92/D gnd DFFSR_192/D vdd OAI22X1
XOAI22X1_81 OAI22X1_81/A OAI22X1_81/B OAI22X1_81/C OAI22X1_81/D gnd OAI22X1_81/Y vdd
+ OAI22X1
XFILL_20_6_0 gnd vdd FILL
XFILL_28_7_0 gnd vdd FILL
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XFILL_3_7_0 gnd vdd FILL
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XFILL_11_6_0 gnd vdd FILL
XCLKBUF1_7 CLKBUF1_7/A gnd CLKBUF1_7/Y vdd CLKBUF1
XNOR2X1_216 INVX8_24/Y NOR2X1_232/B gnd MUX2X1_22/S vdd NOR2X1
XBUFX4_123 DFFSR_245/Q gnd BUFX4_123/Y vdd BUFX4
XBUFX4_167 INVX8_21/Y gnd MUX2X1_26/S vdd BUFX4
XBUFX4_156 INVX8_14/Y gnd BUFX4_156/Y vdd BUFX4
XFILL_19_7_0 gnd vdd FILL
XNOR2X1_238 INVX8_25/Y NOR2X1_238/B gnd MUX2X1_38/S vdd NOR2X1
XBUFX4_134 BUFX4_135/A gnd BUFX4_134/Y vdd BUFX4
XBUFX4_101 AND2X2_1/Y gnd BUFX4_101/Y vdd BUFX4
XNOR2X1_249 INVX8_24/Y NOR2X1_251/B gnd MUX2X1_46/S vdd NOR2X1
XBUFX4_145 INVX8_16/Y gnd BUFX4_145/Y vdd BUFX4
XBUFX4_189 wb_sel_i[2] gnd BUFX4_189/Y vdd BUFX4
XNOR2X1_227 INVX1_156/A BUFX4_157/Y gnd NOR2X1_227/Y vdd NOR2X1
XNOR2X1_205 BUFX4_251/Y INVX1_148/A gnd NOR2X1_205/Y vdd NOR2X1
XBUFX4_112 wb_sel_i[0] gnd MUX2X1_47/S vdd BUFX4
XBUFX4_178 BUFX4_179/A gnd BUFX4_178/Y vdd BUFX4
XINVX8_9 INVX8_9/A gnd OR2X2_1/A vdd INVX8
XBUFX4_18 BUFX4_9/A gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 INVX8_3/Y gnd BUFX4_29/Y vdd BUFX4
XINVX2_156 NOR2X1_19/Y gnd INVX2_156/Y vdd INVX2
XINVX2_101 INVX1_34/A gnd INVX2_101/Y vdd INVX2
XINVX2_112 INVX1_38/A gnd INVX2_112/Y vdd INVX2
XINVX2_123 INVX2_123/A gnd INVX2_123/Y vdd INVX2
XINVX2_145 INVX2_145/A gnd INVX2_145/Y vdd INVX2
XINVX2_134 INVX1_31/A gnd INVX2_134/Y vdd INVX2
XFILL_22_1 gnd vdd FILL
XOAI21X1_508 INVX2_104/Y BUFX4_90/Y OAI21X1_508/C gnd OAI21X1_509/B vdd OAI21X1
XOAI21X1_519 BUFX4_153/Y OAI21X1_519/B OAI21X1_519/C gnd AOI22X1_70/C vdd OAI21X1
XFILL_25_5_0 gnd vdd FILL
XFILL_0_5_0 gnd vdd FILL
XAOI21X1_171 NOR2X1_199/Y BUFX4_154/Y OAI21X1_524/Y gnd OAI22X1_107/C vdd AOI21X1
XAOI21X1_193 INVX2_101/Y OAI21X1_568/B BUFX4_257/Y gnd OAI21X1_568/C vdd AOI21X1
XAOI21X1_182 INVX2_107/Y OAI21X1_547/B INVX8_23/A gnd OAI21X1_547/C vdd AOI21X1
XAOI21X1_160 NOR2X1_182/Y BUFX4_153/Y OAI21X1_495/Y gnd OAI22X1_99/C vdd AOI21X1
XOAI22X1_114 MUX2X1_2/A BUFX4_164/Y OAI22X1_114/C OAI22X1_114/D gnd DFFSR_159/D vdd
+ OAI22X1
XOAI22X1_103 INVX2_90/Y BUFX4_162/Y OAI22X1_103/C OAI22X1_103/D gnd DFFSR_177/D vdd
+ OAI22X1
XFILL_8_6_0 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XNAND3X1_142 NOR3X1_4/B NAND3X1_142/B NAND3X1_142/C gnd NAND3X1_158/B vdd NAND3X1
XNAND3X1_153 MUX2X1_38/B BUFX4_49/Y BUFX4_138/Y gnd NAND3X1_155/B vdd NAND3X1
XNAND3X1_197 BUFX4_65/Y NAND3X1_197/B NAND3X1_197/C gnd AOI21X1_49/B vdd NAND3X1
XNAND3X1_131 INVX2_92/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_133/B vdd NAND3X1
XNAND3X1_175 BUFX4_206/Y NAND3X1_175/B NAND3X1_175/C gnd AOI21X1_46/A vdd NAND3X1
XNAND3X1_164 MUX2X1_18/B BUFX4_47/Y BUFX4_141/Y gnd NAND3X1_166/B vdd NAND3X1
XNAND3X1_186 INVX2_115/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_188/B vdd NAND3X1
XNAND3X1_120 INVX2_76/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_122/B vdd NAND3X1
XOAI21X1_305 BUFX4_178/Y INVX1_94/A BUFX4_34/Y gnd OAI22X1_68/A vdd OAI21X1
XDFFSR_173 INVX2_80/A DFFSR_98/CLK BUFX4_14/Y vdd DFFSR_173/D gnd vdd DFFSR
XDFFSR_151 INVX2_65/A CLKBUF1_20/Y BUFX4_12/Y vdd DFFSR_151/D gnd vdd DFFSR
XBUFX4_3 BUFX4_7/A gnd BUFX4_3/Y vdd BUFX4
XOAI21X1_327 NOR2X1_96/B MUX2X1_41/B BUFX4_39/Y gnd OAI22X1_76/D vdd OAI21X1
XDFFSR_184 INVX1_30/A CLKBUF1_7/Y BUFX4_9/Y vdd DFFSR_184/D gnd vdd DFFSR
XDFFSR_162 INVX1_60/A CLKBUF1_25/Y BUFX4_11/Y vdd DFFSR_162/D gnd vdd DFFSR
XDFFSR_140 MUX2X1_27/B DFFSR_5/CLK BUFX4_11/Y vdd DFFSR_140/D gnd vdd DFFSR
XOAI21X1_338 OAI22X1_79/Y OAI22X1_80/Y NOR2X1_85/Y gnd OAI21X1_338/Y vdd OAI21X1
XOAI21X1_316 BUFX4_179/Y INVX1_99/A BUFX4_36/Y gnd OAI22X1_72/D vdd OAI21X1
XOAI21X1_349 INVX2_68/Y BUFX4_89/Y OAI21X1_672/C gnd AOI21X1_79/B vdd OAI21X1
XDFFSR_195 INVX2_70/A CLKBUF1_54/Y BUFX4_17/Y vdd DFFSR_195/D gnd vdd DFFSR
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 NAND3X1_7/A OAI21X1_7/Y BUFX4_99/Y gnd OAI21X1_8/C vdd NAND3X1
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 AND2X2_3/Y INVX2_35/Y NAND3X1_56/Y gnd DFFSR_59/D vdd OAI21X1
XOAI21X1_124 AND2X2_3/Y INVX2_46/Y NAND3X1_67/Y gnd DFFSR_54/D vdd OAI21X1
XOAI21X1_146 BUFX4_30/Y BUFX4_124/Y INVX1_13/A gnd BUFX2_23/A vdd OAI21X1
XOAI21X1_135 BUFX4_31/Y BUFX4_120/Y INVX2_3/A gnd BUFX2_12/A vdd OAI21X1
XOAI21X1_113 INVX2_41/Y MUX2X1_43/S OAI21X1_81/C gnd NAND3X1_62/B vdd OAI21X1
XOAI21X1_168 XNOR2X1_1/A NOR2X1_42/Y NOR2X1_47/B gnd OAI21X1_169/C vdd OAI21X1
XOAI21X1_179 INVX8_10/Y OR2X2_1/A INVX2_32/A gnd OAI21X1_180/C vdd OAI21X1
XOAI21X1_157 BUFX4_28/Y BUFX4_120/Y INVX1_8/A gnd BUFX2_34/A vdd OAI21X1
XNAND2X1_130 AOI21X1_68/B OAI21X1_236/C gnd XNOR2X1_13/A vdd NAND2X1
XNAND2X1_152 NOR2X1_148/Y NOR2X1_71/Y gnd AOI21X1_84/B vdd NAND2X1
XNAND2X1_185 BUFX4_25/Y wb_dat_i[10] gnd OAI21X1_638/C vdd NAND2X1
XNAND2X1_141 OAI21X1_296/Y OAI21X1_301/Y gnd OAI21X1_302/B vdd NAND2X1
XNAND2X1_163 wb_dat_i[22] MUX2X1_29/S gnd OAI21X1_528/C vdd NAND2X1
XNAND2X1_174 BUFX4_189/Y wb_dat_i[17] gnd OAI21X1_621/C vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_196 MUX2X1_35/S wb_dat_i[4] gnd OAI21X1_651/C vdd NAND2X1
XFILL_13_3_0 gnd vdd FILL
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XAOI22X1_19 INVX8_6/Y INVX2_80/A INVX2_82/A INVX8_7/Y gnd NAND3X1_81/C vdd AOI22X1
XOAI21X1_691 INVX2_77/Y MUX2X1_37/S OAI21X1_693/C gnd OAI21X1_691/Y vdd OAI21X1
XOAI21X1_680 NOR2X1_248/Y INVX2_78/Y BUFX4_234/Y gnd OAI21X1_680/Y vdd OAI21X1
XBUFX2_51 DFFSR_80/Q gnd wb_dat_o[15] vdd BUFX2
XBUFX2_40 DFFSR_69/Q gnd wb_dat_o[4] vdd BUFX2
XBUFX2_62 DFFSR_91/Q gnd wb_dat_o[26] vdd BUFX2
XBUFX2_73 INVX4_6/A gnd BUFX2_73/Y vdd BUFX2
XAOI21X1_52 AOI21X1_52/A AOI21X1_52/B INVX8_13/Y gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_41 AOI21X1_41/A AOI21X1_41/B INVX2_66/Y gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_30 NAND2X1_97/Y NAND2X1_99/Y INVX2_55/A gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_74 INVX4_7/A INVX4_8/A BUFX4_272/Y gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_63 AOI21X1_63/A AOI21X1_63/B INVX4_3/A gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_85 BUFX4_264/Y AOI21X1_85/B BUFX4_250/Y gnd AOI22X1_38/D vdd AOI21X1
XOAI21X1_3 INVX1_2/Y BUFX4_89/Y OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XAOI21X1_96 INVX2_97/Y AOI21X1_96/B BUFX4_268/Y gnd AOI21X1_96/Y vdd AOI21X1
XOAI22X1_93 MUX2X1_5/A BUFX4_43/Y OAI22X1_93/C OAI22X1_93/D gnd DFFSR_191/D vdd OAI22X1
XOAI22X1_82 OAI22X1_82/A OAI22X1_82/B OAI22X1_82/C OAI22X1_82/D gnd OAI22X1_82/Y vdd
+ OAI22X1
XOAI22X1_60 OAI22X1_60/A NOR2X1_97/Y NOR2X1_98/Y OAI22X1_60/D gnd OAI22X1_60/Y vdd
+ OAI22X1
XOAI22X1_71 OAI22X1_71/A OAI22X1_71/B OAI22X1_71/C OAI22X1_71/D gnd OAI22X1_71/Y vdd
+ OAI22X1
XFILL_20_6_1 gnd vdd FILL
XFILL_28_7_1 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XXOR2X1_6 OR2X2_8/A XOR2X1_6/B gnd XOR2X1_6/Y vdd XOR2X1
XFILL_2_2_0 gnd vdd FILL
XFILL_3_7_1 gnd vdd FILL
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_9/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_11_6_1 gnd vdd FILL
XCLKBUF1_8 CLKBUF1_8/A gnd DFFSR_4/CLK vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XBUFX4_102 AND2X2_1/Y gnd BUFX4_102/Y vdd BUFX4
XNOR2X1_217 INVX8_24/Y NOR2X1_233/B gnd AND2X2_21/B vdd NOR2X1
XFILL_19_7_1 gnd vdd FILL
XBUFX4_168 NOR3X1_9/Y gnd BUFX4_168/Y vdd BUFX4
XFILL_18_2_0 gnd vdd FILL
XBUFX4_146 INVX8_16/Y gnd BUFX4_146/Y vdd BUFX4
XBUFX4_157 INVX8_14/Y gnd BUFX4_157/Y vdd BUFX4
XNOR2X1_228 INVX8_24/Y NOR2X1_243/B gnd NOR2X1_228/Y vdd NOR2X1
XNOR2X1_239 INVX8_25/Y NOR2X1_239/B gnd NOR2X1_239/Y vdd NOR2X1
XBUFX4_113 BUFX4_117/A gnd BUFX4_113/Y vdd BUFX4
XBUFX4_124 DFFSR_245/Q gnd BUFX4_124/Y vdd BUFX4
XBUFX4_179 BUFX4_179/A gnd BUFX4_179/Y vdd BUFX4
XNOR2X1_206 BUFX4_179/Y INVX1_138/Y gnd INVX4_12/A vdd NOR2X1
XBUFX4_135 BUFX4_135/A gnd OAI22X1_7/D vdd BUFX4
XBUFX4_19 wb_sel_i[1] gnd BUFX4_19/Y vdd BUFX4
XINVX2_102 INVX1_33/A gnd INVX2_102/Y vdd INVX2
XINVX2_157 INVX2_157/A gnd INVX2_157/Y vdd INVX2
XINVX2_146 NOR2X1_96/A gnd INVX2_146/Y vdd INVX2
XINVX2_135 INVX1_30/A gnd INVX2_135/Y vdd INVX2
XINVX2_113 INVX1_37/A gnd INVX2_113/Y vdd INVX2
XINVX2_124 INVX1_26/A gnd INVX2_124/Y vdd INVX2
XOAI21X1_509 BUFX4_150/Y OAI21X1_509/B BUFX4_165/Y gnd OAI22X1_102/D vdd OAI21X1
XFILL_25_5_1 gnd vdd FILL
XFILL_0_5_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 INVX2_108/Y OAI21X1_465/B BUFX4_254/Y gnd OAI21X1_465/C vdd AOI21X1
XAOI21X1_194 BUFX4_257/Y OAI21X1_569/Y BUFX4_4/Y gnd AOI22X1_77/D vdd AOI21X1
XAOI21X1_172 AND2X2_18/Y BUFX4_157/Y OAI21X1_527/Y gnd OAI22X1_108/C vdd AOI21X1
XAOI21X1_161 NOR2X1_183/Y BUFX4_155/Y OAI21X1_498/Y gnd OAI22X1_100/C vdd AOI21X1
XAOI21X1_183 BUFX4_259/Y OAI21X1_548/Y BUFX4_5/Y gnd AOI22X1_74/D vdd AOI21X1
XOAI22X1_115 MUX2X1_6/A BUFX4_164/Y OAI22X1_115/C OAI22X1_115/D gnd DFFSR_157/D vdd
+ OAI22X1
XOAI22X1_104 MUX2X1_15/B MUX2X1_26/S OAI22X1_104/C OAI22X1_104/D gnd DFFSR_176/D vdd
+ OAI22X1
XFILL_7_1_0 gnd vdd FILL
XFILL_8_6_1 gnd vdd FILL
XNAND3X1_121 INVX2_77/Y BUFX4_50/Y BUFX4_137/Y gnd NAND3X1_122/C vdd NAND3X1
XNAND3X1_110 INVX2_70/Y BUFX4_75/Y BUFX4_58/Y gnd AOI21X1_37/B vdd NAND3X1
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XNAND3X1_132 INVX2_93/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_133/C vdd NAND3X1
XNAND3X1_154 INVX2_102/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_155/C vdd NAND3X1
XNAND3X1_187 INVX2_116/Y BUFX4_48/Y BUFX4_137/Y gnd NAND3X1_188/C vdd NAND3X1
XNAND3X1_198 INVX2_121/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_200/B vdd NAND3X1
XNAND3X1_176 MUX2X1_30/B BUFX4_46/Y BUFX4_141/Y gnd NAND3X1_178/B vdd NAND3X1
XNAND3X1_165 INVX2_105/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_166/C vdd NAND3X1
XNAND3X1_143 INVX2_97/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_145/B vdd NAND3X1
XOAI21X1_328 OAI22X1_75/Y OAI22X1_76/Y INVX2_154/Y gnd OAI21X1_328/Y vdd OAI21X1
XOAI21X1_317 OAI22X1_71/Y OAI22X1_72/Y NOR2X1_85/Y gnd OAI21X1_317/Y vdd OAI21X1
XOAI21X1_306 BUFX4_178/Y INVX1_95/A BUFX4_36/Y gnd OAI22X1_68/D vdd OAI21X1
XDFFSR_141 MUX2X1_25/B CLKBUF1_49/Y BUFX4_14/Y vdd MUX2X1_26/Y gnd vdd DFFSR
XDFFSR_185 INVX1_33/A CLKBUF1_2/Y BUFX4_18/Y vdd DFFSR_185/D gnd vdd DFFSR
XDFFSR_163 INVX2_71/A CLKBUF1_21/Y BUFX4_10/Y vdd DFFSR_163/D gnd vdd DFFSR
XBUFX4_4 BUFX4_7/A gnd BUFX4_4/Y vdd BUFX4
XDFFSR_130 MUX2X1_31/B CLKBUF1_35/Y BUFX4_11/Y vdd DFFSR_130/D gnd vdd DFFSR
XDFFSR_196 NOR2X1_98/A CLKBUF1_20/Y BUFX4_9/Y vdd DFFSR_196/D gnd vdd DFFSR
XDFFSR_152 INVX1_31/A CLKBUF1_15/Y BUFX4_11/Y vdd DFFSR_152/D gnd vdd DFFSR
XOAI21X1_339 INVX2_115/A NOR2X1_89/B BUFX4_78/Y gnd OAI22X1_81/D vdd OAI21X1
XDFFSR_174 INVX2_116/A CLKBUF1_40/Y BUFX4_10/Y vdd DFFSR_174/D gnd vdd DFFSR
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 NAND3X1_7/A OAI21X1_9/Y BUFX4_99/Y gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_169 INVX1_69/Y NOR2X1_47/B OAI21X1_169/C gnd DFFSR_104/D vdd OAI21X1
XOAI21X1_158 OR2X2_2/Y NAND2X1_77/Y INVX8_9/A gnd NOR2X1_46/B vdd OAI21X1
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_103 INVX2_36/Y BUFX4_22/Y OAI21X1_73/C gnd NAND3X1_57/B vdd OAI21X1
XOAI21X1_136 BUFX4_27/Y INVX8_9/A INVX2_4/A gnd BUFX2_13/A vdd OAI21X1
XOAI21X1_125 INVX4_1/Y NAND2X1_34/Y NOR2X1_17/B gnd BUFX4_117/A vdd OAI21X1
XOAI21X1_147 BUFX4_30/Y BUFX4_120/Y INVX1_14/A gnd BUFX2_24/A vdd OAI21X1
XOAI21X1_114 AND2X2_3/Y INVX2_41/Y NAND3X1_62/Y gnd DFFSR_49/D vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd mosi_pad_o vdd BUFX2
XNAND2X1_120 INVX2_151/A AND2X2_12/B gnd NOR3X1_7/C vdd NAND2X1
XNAND2X1_131 BUFX2_80/A XNOR2X1_13/Y gnd NAND2X1_132/B vdd NAND2X1
XNAND2X1_153 BUFX4_87/Y wb_dat_i[28] gnd OAI21X1_514/C vdd NAND2X1
XNAND2X1_164 NOR2X1_71/Y NOR2X1_154/Y gnd AOI21X1_96/B vdd NAND2X1
XNAND2X1_142 OAI21X1_307/Y OAI21X1_312/Y gnd OAI21X1_323/A vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_175 NOR2X1_160/Y NOR2X1_71/Y gnd OAI21X1_377/B vdd NAND2X1
XNAND2X1_197 NOR2X1_156/Y INVX1_139/A gnd OAI21X1_401/B vdd NAND2X1
XNAND2X1_186 INVX1_143/A INVX8_14/A gnd NAND2X1_186/Y vdd NAND2X1
XINVX2_1 wb_adr_i[2] gnd INVX2_1/Y vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XAOI21X1_1 MUX2X1_43/B BUFX4_115/Y OAI22X1_3/Y gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_670 INVX2_73/Y BUFX4_187/Y OAI21X1_697/C gnd OAI21X1_670/Y vdd OAI21X1
XOAI21X1_681 INVX2_78/Y MUX2X1_35/S OAI21X1_693/C gnd OAI21X1_682/B vdd OAI21X1
XOAI21X1_692 BUFX4_160/Y OAI21X1_692/B OAI21X1_692/C gnd AOI22X1_89/C vdd OAI21X1
XBUFX2_41 DFFSR_70/Q gnd wb_dat_o[5] vdd BUFX2
XBUFX2_74 INVX2_52/A gnd BUFX2_74/Y vdd BUFX2
XBUFX2_30 BUFX2_30/A gnd ss_pad_o[27] vdd BUFX2
XBUFX2_52 DFFSR_81/Q gnd wb_dat_o[16] vdd BUFX2
XBUFX2_63 DFFSR_92/Q gnd wb_dat_o[27] vdd BUFX2
XAOI21X1_75 INVX1_131/Y AOI21X1_75/B NOR2X1_73/B gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_64 INVX2_48/A NOR3X1_5/Y OR2X2_4/B gnd NOR3X1_6/B vdd AOI21X1
XAOI21X1_20 NOR2X1_28/A AND2X2_6/A AND2X2_5/Y gnd AOI21X1_20/Y vdd AOI21X1
XAOI21X1_42 AOI21X1_42/A AOI21X1_42/B INVX2_55/Y gnd NOR3X1_4/C vdd AOI21X1
XAOI21X1_31 AOI21X1_31/A AOI21X1_31/B INVX2_55/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_86 MUX2X1_4/B AOI21X1_86/B BUFX4_263/Y gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_53 AOI21X1_53/A AOI21X1_53/B BUFX4_81/Y gnd AOI21X1_53/Y vdd AOI21X1
XOAI21X1_4 OAI21X1_8/A INVX1_2/Y OAI21X1_4/C gnd DFFSR_26/D vdd OAI21X1
XAOI21X1_97 BUFX4_265/Y AOI21X1_97/B BUFX4_246/Y gnd AOI22X1_44/D vdd AOI21X1
XOAI22X1_50 INVX1_66/Y NOR2X1_47/B OAI22X1_50/C INVX1_79/Y gnd DFFSR_115/D vdd OAI22X1
XOAI22X1_61 OAI22X1_61/A NOR2X1_99/Y OAI22X1_61/C OAI22X1_61/D gnd OAI22X1_61/Y vdd
+ OAI22X1
XOAI22X1_83 INVX2_88/Y BUFX4_43/Y OAI22X1_83/C OAI22X1_83/D gnd DFFSR_209/D vdd OAI22X1
XOAI22X1_94 INVX2_120/Y BUFX4_41/Y OAI22X1_94/C OAI22X1_94/D gnd DFFSR_190/D vdd OAI22X1
XOAI22X1_72 OAI22X1_72/A OAI22X1_72/B OAI22X1_72/C OAI22X1_72/D gnd OAI22X1_72/Y vdd
+ OAI22X1
XFILL_3_1 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A MUX2X1_8/B MUX2X1_8/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 CLKBUF1_9/A gnd CLKBUF1_9/Y vdd CLKBUF1
XBUFX4_136 BUFX4_142/A gnd BUFX4_136/Y vdd BUFX4
XBUFX4_125 DFFSR_245/Q gnd BUFX4_125/Y vdd BUFX4
XBUFX4_103 AND2X2_1/Y gnd OAI21X1_8/A vdd BUFX4
XBUFX4_114 BUFX4_117/A gnd BUFX4_114/Y vdd BUFX4
XNOR2X1_207 INVX4_12/Y INVX1_150/Y gnd NOR2X1_207/Y vdd NOR2X1
XBUFX4_147 INVX8_23/Y gnd BUFX4_147/Y vdd BUFX4
XFILL_18_2_1 gnd vdd FILL
XBUFX4_158 INVX8_14/Y gnd BUFX4_158/Y vdd BUFX4
XBUFX4_169 NOR3X1_9/Y gnd BUFX4_169/Y vdd BUFX4
XNOR2X1_229 BUFX4_179/Y INVX1_149/Y gnd INVX8_25/A vdd NOR2X1
XNOR2X1_218 INVX8_24/Y NOR2X1_234/B gnd MUX2X1_24/S vdd NOR2X1
XINVX2_103 INVX2_103/A gnd INVX2_103/Y vdd INVX2
XINVX2_114 INVX1_36/A gnd INVX2_114/Y vdd INVX2
XINVX2_158 NOR2X1_94/Y gnd INVX2_158/Y vdd INVX2
XINVX2_147 NOR2X1_98/A gnd INVX2_147/Y vdd INVX2
XINVX2_136 INVX2_136/A gnd INVX2_136/Y vdd INVX2
XINVX2_125 INVX1_25/A gnd INVX2_125/Y vdd INVX2
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_184 NOR2X1_207/Y BUFX4_154/Y OAI21X1_549/Y gnd OAI22X1_112/C vdd AOI21X1
XAOI21X1_151 NOR2X1_174/Y BUFX4_154/Y OAI21X1_468/Y gnd OAI22X1_91/C vdd AOI21X1
XAOI21X1_162 NOR2X1_184/Y BUFX4_153/Y OAI21X1_501/Y gnd OAI22X1_101/C vdd AOI21X1
XAOI21X1_140 NOR2X1_168/Y BUFX4_160/Y OAI21X1_426/Y gnd OAI22X1_86/C vdd AOI21X1
XAOI21X1_173 AND2X2_19/Y BUFX4_159/Y OAI21X1_530/Y gnd OAI22X1_109/C vdd AOI21X1
XAOI21X1_195 INVX2_134/Y OAI21X1_570/B INVX8_23/A gnd OAI21X1_570/C vdd AOI21X1
XOAI22X1_105 MUX2X1_2/B BUFX4_164/Y OAI22X1_105/C OAI22X1_105/D gnd DFFSR_175/D vdd
+ OAI22X1
XOAI22X1_116 INVX2_143/Y BUFX4_162/Y OAI22X1_116/C OAI22X1_116/D gnd DFFSR_156/D vdd
+ OAI22X1
XFILL_7_1_1 gnd vdd FILL
XNAND3X1_155 BUFX4_63/Y NAND3X1_155/B NAND3X1_155/C gnd NAND3X1_156/C vdd NAND3X1
XNAND3X1_111 INVX2_71/Y BUFX4_48/Y BUFX4_138/Y gnd AOI21X1_38/A vdd NAND3X1
XFILL_15_0_1 gnd vdd FILL
XNAND3X1_133 BUFX4_204/Y NAND3X1_133/B NAND3X1_133/C gnd NAND3X1_134/C vdd NAND3X1
XNAND3X1_144 INVX2_98/Y BUFX4_47/Y BUFX4_141/Y gnd NAND3X1_145/C vdd NAND3X1
XNAND3X1_166 BUFX4_64/Y NAND3X1_166/B NAND3X1_166/C gnd AOI21X1_44/B vdd NAND3X1
XNAND3X1_100 BUFX4_65/Y NAND3X1_98/Y NAND3X1_99/Y gnd AOI21X1_34/A vdd NAND3X1
XNAND3X1_122 BUFX4_205/Y NAND3X1_122/B NAND3X1_122/C gnd AOI21X1_40/A vdd NAND3X1
XNAND3X1_188 BUFX4_205/Y NAND3X1_188/B NAND3X1_188/C gnd AOI21X1_48/A vdd NAND3X1
XNAND3X1_199 INVX2_122/Y BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_200/C vdd NAND3X1
XNAND3X1_177 INVX2_111/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_178/C vdd NAND3X1
XOAI21X1_318 INVX2_57/A NOR2X1_84/B BUFX4_77/Y gnd OAI22X1_73/D vdd OAI21X1
XOAI21X1_329 INVX2_103/A BUFX4_222/Y BUFX4_79/Y gnd OAI22X1_77/D vdd OAI21X1
XOAI21X1_307 OAI22X1_67/Y OAI22X1_68/Y INVX2_154/Y gnd OAI21X1_307/Y vdd OAI21X1
XDFFSR_175 INVX2_54/A DFFSR_70/CLK BUFX4_14/Y vdd DFFSR_175/D gnd vdd DFFSR
XDFFSR_153 INVX1_34/A CLKBUF1_9/Y BUFX4_10/Y vdd DFFSR_153/D gnd vdd DFFSR
XDFFSR_131 INVX1_97/A DFFSR_86/CLK BUFX4_11/Y vdd DFFSR_131/D gnd vdd DFFSR
XDFFSR_197 INVX2_91/A CLKBUF1_16/Y BUFX4_12/Y vdd DFFSR_197/D gnd vdd DFFSR
XDFFSR_164 NOR2X1_96/A CLKBUF1_6/A BUFX4_12/Y vdd DFFSR_164/D gnd vdd DFFSR
XDFFSR_120 INVX1_118/A CLKBUF1_6/A BUFX4_13/Y vdd DFFSR_120/D gnd vdd DFFSR
XDFFSR_142 MUX2X1_23/B DFFSR_82/CLK BUFX4_11/Y vdd DFFSR_142/D gnd vdd DFFSR
XBUFX4_5 BUFX4_7/A gnd BUFX4_5/Y vdd BUFX4
XDFFSR_186 INVX1_36/A CLKBUF1_49/Y BUFX4_10/Y vdd DFFSR_186/D gnd vdd DFFSR
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XNAND3X1_8 AND2X2_1/B NAND3X1_8/B BUFX4_95/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_159 INVX8_10/Y OR2X2_1/A INVX2_39/A gnd OAI21X1_160/C vdd OAI21X1
XOAI21X1_115 INVX2_42/Y BUFX4_108/Y OAI21X1_83/C gnd NAND3X1_63/B vdd OAI21X1
XOAI21X1_104 AND2X2_3/Y INVX2_36/Y NAND3X1_57/Y gnd DFFSR_60/D vdd OAI21X1
XOAI21X1_126 BUFX4_29/Y BUFX4_118/Y DFFSR_1/Q gnd BUFX2_3/A vdd OAI21X1
XOAI21X1_148 BUFX4_30/Y BUFX4_124/Y INVX1_15/A gnd BUFX2_25/A vdd OAI21X1
XOAI21X1_137 BUFX4_28/Y BUFX4_120/Y INVX2_5/A gnd BUFX2_14/A vdd OAI21X1
XBUFX2_2 OR2X2_1/B gnd sclk_pad_o vdd BUFX2
XNAND2X1_121 INVX1_128/A AOI21X1_66/Y gnd AOI22X1_34/D vdd NAND2X1
XNAND2X1_132 NAND2X1_132/A NAND2X1_132/B gnd NOR2X1_94/B vdd NAND2X1
XNAND2X1_110 MUX2X1_15/Y NOR2X1_66/B gnd NAND3X1_213/A vdd NAND2X1
XNAND2X1_143 OAI21X1_317/Y OAI21X1_322/Y gnd OAI21X1_323/B vdd NAND2X1
XNAND2X1_187 NOR2X1_151/Y INVX1_139/A gnd OAI21X1_391/B vdd NAND2X1
XNAND2X1_154 NOR2X1_149/Y NOR2X1_71/Y gnd AOI21X1_86/B vdd NAND2X1
XNAND2X1_165 BUFX4_188/Y wb_dat_i[21] gnd OAI21X1_605/C vdd NAND2X1
XNAND2X1_176 NAND2X1_9/B wb_dat_i[16] gnd OAI21X1_624/C vdd NAND2X1
XNAND2X1_198 BUFX4_111/Y wb_dat_i[3] gnd OAI21X1_573/C vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_660 NOR2X1_242/Y OAI21X1_660/B OAI21X1_660/C gnd DFFSR_117/D vdd OAI21X1
XAOI21X1_2 INVX1_104/A BUFX4_115/Y OAI22X1_6/Y gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_671 BUFX4_153/Y OAI21X1_671/B OAI21X1_671/C gnd AOI22X1_84/C vdd OAI21X1
XOAI21X1_682 BUFX4_234/Y OAI21X1_682/B BUFX4_45/Y gnd OAI22X1_120/D vdd OAI21X1
XOAI21X1_693 INVX2_76/Y BUFX4_111/Y OAI21X1_693/C gnd OAI21X1_693/Y vdd OAI21X1
XXNOR2X1_10 INVX1_126/A XOR2X1_3/Y gnd INVX1_128/A vdd XNOR2X1
XBUFX2_64 DFFSR_93/Q gnd wb_dat_o[28] vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd ss_pad_o[28] vdd BUFX2
XBUFX2_75 NOR3X1_6/A gnd BUFX2_75/Y vdd BUFX2
XBUFX2_53 DFFSR_82/Q gnd wb_dat_o[17] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd ss_pad_o[17] vdd BUFX2
XBUFX2_42 DFFSR_71/Q gnd wb_dat_o[6] vdd BUFX2
XFILL_23_6_0 gnd vdd FILL
XAOI21X1_65 INVX1_126/A INVX1_125/Y INVX2_51/Y gnd NOR3X1_7/B vdd AOI21X1
XAOI21X1_21 NOR2X1_43/B NOR2X1_25/Y OR2X2_1/A gnd NOR2X1_47/B vdd AOI21X1
XAOI21X1_76 INVX1_134/Y AOI21X1_77/B NOR3X1_9/B gnd BUFX4_39/A vdd AOI21X1
XAOI21X1_10 INVX1_100/A BUFX4_117/Y OAI22X1_30/Y gnd NAND2X1_44/A vdd AOI21X1
XAOI21X1_43 AOI21X1_43/A AOI21X1_43/B INVX2_55/A gnd NOR3X1_4/A vdd AOI21X1
XAOI21X1_87 BUFX4_263/Y AOI21X1_87/B BUFX4_243/Y gnd AOI22X1_39/D vdd AOI21X1
XAOI21X1_32 NAND2X1_92/A NAND3X1_91/Y XOR2X1_3/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_54 AOI21X1_54/A AOI21X1_54/B NOR3X1_4/B gnd AOI21X1_54/Y vdd AOI21X1
XOAI21X1_5 INVX1_3/Y BUFX4_91/Y OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_98 INVX2_136/Y AOI21X1_98/B BUFX4_266/Y gnd AOI21X1_98/Y vdd AOI21X1
XFILL_6_7_0 gnd vdd FILL
XFILL_14_6_0 gnd vdd FILL
XOAI22X1_95 MUX2X1_7/A BUFX4_44/Y OAI22X1_95/C OAI22X1_95/D gnd DFFSR_189/D vdd OAI22X1
XOAI22X1_84 MUX2X1_14/B BUFX4_44/Y OAI22X1_84/C OAI22X1_84/D gnd DFFSR_208/D vdd OAI22X1
XOAI22X1_62 OAI22X1_62/A OAI22X1_62/B OAI22X1_62/C OAI22X1_62/D gnd OAI22X1_62/Y vdd
+ OAI22X1
XOAI22X1_73 OAI22X1_73/A OAI22X1_73/B OAI22X1_73/C OAI22X1_73/D gnd OAI22X1_73/Y vdd
+ OAI22X1
XOAI22X1_40 OAI22X1_5/A INVX2_7/Y INVX2_36/Y OAI22X1_5/D gnd NOR2X1_15/A vdd OAI22X1
XOAI22X1_51 OAI22X1_51/A NOR2X1_77/Y NOR2X1_78/Y OAI22X1_51/D gnd OAI22X1_51/Y vdd
+ OAI22X1
XOAI21X1_490 INVX2_102/Y MUX2X1_47/S OAI21X1_569/C gnd OAI21X1_491/B vdd OAI21X1
XFILL_3_2 gnd vdd FILL
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XBUFX4_148 INVX8_23/Y gnd BUFX4_148/Y vdd BUFX4
XBUFX4_115 BUFX4_117/A gnd BUFX4_115/Y vdd BUFX4
XBUFX4_104 AND2X2_1/Y gnd OAI21X1_6/A vdd BUFX4
XBUFX4_159 INVX8_14/Y gnd BUFX4_159/Y vdd BUFX4
XBUFX4_126 DFFSR_245/Q gnd BUFX4_126/Y vdd BUFX4
XBUFX4_137 BUFX4_142/A gnd BUFX4_137/Y vdd BUFX4
XNOR2X1_208 INVX4_12/Y INVX1_151/Y gnd NOR2X1_208/Y vdd NOR2X1
XNOR2X1_219 INVX8_24/Y NOR2X1_235/B gnd NOR2X1_219/Y vdd NOR2X1
XFILL_20_4_0 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XFILL_3_5_0 gnd vdd FILL
XINVX2_137 INVX2_137/A gnd INVX2_137/Y vdd INVX2
XINVX2_104 INVX2_104/A gnd INVX2_104/Y vdd INVX2
XINVX2_126 INVX1_24/A gnd INVX2_126/Y vdd INVX2
XINVX2_115 INVX2_115/A gnd INVX2_115/Y vdd INVX2
XFILL_11_4_0 gnd vdd FILL
XINVX2_159 INVX2_159/A gnd INVX2_159/Y vdd INVX2
XINVX2_148 INVX1_20/A gnd INVX2_148/Y vdd INVX2
XFILL_19_5_0 gnd vdd FILL
XAOI21X1_185 NOR2X1_208/Y BUFX4_152/Y OAI21X1_552/Y gnd OAI22X1_113/C vdd AOI21X1
XAOI21X1_141 NOR2X1_169/Y BUFX4_152/Y OAI21X1_430/Y gnd OAI22X1_87/C vdd AOI21X1
XAOI21X1_152 NOR2X1_175/Y BUFX4_152/Y OAI21X1_471/Y gnd OAI22X1_92/C vdd AOI21X1
XAOI21X1_174 INVX2_137/Y OAI21X1_534/B BUFX4_258/Y gnd OAI21X1_534/C vdd AOI21X1
XAOI21X1_163 INVX2_150/Y OAI21X1_504/B BUFX4_254/Y gnd OAI21X1_504/C vdd AOI21X1
XAOI21X1_196 INVX8_23/A OAI21X1_571/Y BUFX4_7/Y gnd AOI22X1_78/D vdd AOI21X1
XAOI21X1_130 INVX2_124/Y OAI21X1_403/B BUFX4_261/Y gnd OAI21X1_403/C vdd AOI21X1
XOAI22X1_106 MUX2X1_6/B BUFX4_164/Y OAI22X1_106/C OAI22X1_106/D gnd DFFSR_173/D vdd
+ OAI22X1
XOAI22X1_117 INVX2_95/Y BUFX4_166/Y OAI22X1_117/C OAI22X1_117/D gnd DFFSR_149/D vdd
+ OAI22X1
XNAND3X1_156 MUX2X1_9/S NAND3X1_156/B NAND3X1_156/C gnd NAND3X1_157/C vdd NAND3X1
XNAND3X1_112 INVX2_72/Y BUFX4_75/Y BUFX4_58/Y gnd AOI21X1_38/B vdd NAND3X1
XNAND3X1_189 MUX2X1_24/B BUFX4_48/Y BUFX4_137/Y gnd NAND3X1_191/B vdd NAND3X1
XNAND3X1_178 BUFX4_62/Y NAND3X1_178/B NAND3X1_178/C gnd AOI21X1_46/B vdd NAND3X1
XNAND3X1_134 INVX8_13/Y NAND3X1_134/B NAND3X1_134/C gnd NAND3X1_142/B vdd NAND3X1
XNAND3X1_145 BUFX4_206/Y NAND3X1_145/B NAND3X1_145/C gnd NAND3X1_149/B vdd NAND3X1
XNAND3X1_101 INVX2_64/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_103/B vdd NAND3X1
XNAND3X1_123 INVX1_99/Y BUFX4_50/Y BUFX4_136/Y gnd NAND3X1_125/B vdd NAND3X1
XNAND3X1_167 INVX2_106/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_169/B vdd NAND3X1
XFILL_20_1 gnd vdd FILL
XDFFSR_110 INVX1_74/A CLKBUF1_3/Y vdd DFFSR_113/S DFFSR_110/D gnd vdd DFFSR
XDFFSR_143 INVX1_93/A CLKBUF1_41/Y BUFX4_18/Y vdd DFFSR_143/D gnd vdd DFFSR
XOAI21X1_319 INVX2_56/A NOR2X1_84/B BUFX4_168/Y gnd OAI22X1_73/A vdd OAI21X1
XDFFSR_121 MUX2X1_37/B DFFSR_1/CLK BUFX4_18/Y vdd DFFSR_121/D gnd vdd DFFSR
XDFFSR_132 INVX1_122/A CLKBUF1_25/Y BUFX4_13/Y vdd DFFSR_132/D gnd vdd DFFSR
XOAI21X1_308 INVX2_68/A NOR2X1_89/B BUFX4_78/Y gnd OAI22X1_69/D vdd OAI21X1
XDFFSR_176 INVX2_132/A DFFSR_41/CLK BUFX4_14/Y vdd DFFSR_176/D gnd vdd DFFSR
XBUFX4_6 BUFX4_7/A gnd BUFX4_6/Y vdd BUFX4
XDFFSR_198 INVX2_123/A CLKBUF1_10/Y BUFX4_9/Y vdd DFFSR_198/D gnd vdd DFFSR
XDFFSR_165 INVX2_93/A CLKBUF1_6/A BUFX4_13/Y vdd DFFSR_165/D gnd vdd DFFSR
XDFFSR_154 INVX1_37/A CLKBUF1_6/Y BUFX4_11/Y vdd DFFSR_154/D gnd vdd DFFSR
XDFFSR_187 INVX2_78/A CLKBUF1_45/Y BUFX4_10/Y vdd DFFSR_187/D gnd vdd DFFSR
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XFILL_25_3_0 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XNAND3X1_9 NAND3X1_9/A NAND3X1_9/B BUFX4_98/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_116 AND2X2_3/Y INVX2_42/Y NAND3X1_63/Y gnd DFFSR_50/D vdd OAI21X1
XOAI21X1_138 BUFX4_29/Y INVX8_9/A INVX2_6/A gnd BUFX2_15/A vdd OAI21X1
XOAI21X1_127 BUFX4_27/Y INVX8_9/A DFFSR_2/Q gnd BUFX2_4/A vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd ss_pad_o[0] vdd BUFX2
XOAI21X1_149 BUFX4_30/Y BUFX4_124/Y INVX1_16/A gnd BUFX2_26/A vdd OAI21X1
XOAI21X1_105 INVX2_37/Y BUFX4_23/Y OAI21X1_45/C gnd NAND3X1_58/B vdd OAI21X1
XNAND2X1_122 INVX1_127/Y INVX4_8/Y gnd AOI21X1_67/A vdd NAND2X1
XNAND2X1_111 MUX2X1_16/Y BUFX4_66/Y gnd NAND3X1_213/B vdd NAND2X1
XNAND2X1_100 MUX2X1_4/Y NOR2X1_66/B gnd AOI21X1_31/A vdd NAND2X1
XNAND2X1_155 BUFX4_89/Y wb_dat_i[27] gnd OAI21X1_590/C vdd NAND2X1
XNAND2X1_133 NOR2X1_75/Y NOR2X1_71/Y gnd AOI21X1_78/B vdd NAND2X1
XNAND2X1_177 wb_dat_i[14] BUFX4_25/Y gnd OAI21X1_548/C vdd NAND2X1
XNAND2X1_166 NOR2X1_71/Y NOR2X1_155/Y gnd AOI21X1_98/B vdd NAND2X1
XNAND2X1_144 OAI21X1_328/Y OAI21X1_333/Y gnd OAI21X1_344/A vdd NAND2X1
XNAND2X1_188 BUFX4_19/Y wb_dat_i[9] gnd OAI21X1_641/C vdd NAND2X1
XNAND2X1_199 NOR2X1_157/Y INVX1_139/A gnd OAI21X1_403/B vdd NAND2X1
XOAI21X1_650 BUFX4_163/Y MUX2X1_37/Y OAI21X1_650/C gnd DFFSR_121/D vdd OAI21X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_694 INVX1_97/Y BUFX4_24/Y OAI21X1_694/C gnd OAI21X1_694/Y vdd OAI21X1
XOAI21X1_672 INVX2_69/Y BUFX4_91/Y OAI21X1_672/C gnd OAI21X1_672/Y vdd OAI21X1
XOAI21X1_683 BUFX4_121/Y INVX8_22/Y NOR2X1_246/Y gnd NOR2X1_251/B vdd OAI21X1
XAOI21X1_3 MUX2X1_41/B BUFX4_113/Y OAI22X1_9/Y gnd AOI21X1_3/Y vdd AOI21X1
XOAI21X1_661 BUFX4_121/Y INVX8_20/Y MUX2X1_44/Y gnd OAI21X1_662/C vdd OAI21X1
XXNOR2X1_11 XNOR2X1_9/A INVX4_4/Y gnd XNOR2X1_11/Y vdd XNOR2X1
XINVX1_90 XOR2X1_3/Y gnd INVX1_90/Y vdd INVX1
XBUFX2_10 BUFX2_10/A gnd ss_pad_o[7] vdd BUFX2
XBUFX2_76 XOR2X1_3/B gnd BUFX2_76/Y vdd BUFX2
XBUFX2_65 DFFSR_94/Q gnd wb_dat_o[29] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd ss_pad_o[29] vdd BUFX2
XBUFX2_54 DFFSR_83/Q gnd wb_dat_o[18] vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd ss_pad_o[18] vdd BUFX2
XBUFX2_43 DFFSR_72/Q gnd wb_dat_o[7] vdd BUFX2
XNOR2X1_1 INVX8_9/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XFILL_23_6_1 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_66 AOI21X1_66/A NOR3X1_7/Y AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_22 NOR2X1_26/B AND2X2_7/B NOR2X1_43/B gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_77 INVX1_134/Y AOI21X1_77/B NOR3X1_8/A gnd BUFX4_35/A vdd AOI21X1
XAOI21X1_55 AOI21X1_55/A AOI21X1_55/B INVX8_13/A gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_11 INVX1_113/A BUFX4_114/Y OAI22X1_33/Y gnd NAND2X1_45/A vdd AOI21X1
XOAI21X1_6 OAI21X1_6/A INVX1_3/Y OAI21X1_6/C gnd DFFSR_27/D vdd OAI21X1
XAOI21X1_99 BUFX4_266/Y AOI21X1_99/B BUFX4_244/Y gnd AOI22X1_45/D vdd AOI21X1
XAOI21X1_44 AOI21X1_44/A AOI21X1_44/B BUFX4_81/Y gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_33 NAND3X1_94/Y NAND3X1_97/Y INVX8_13/A gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_88 INVX2_115/Y AOI21X1_88/B BUFX4_265/Y gnd AOI21X1_88/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_6_7_1 gnd vdd FILL
XOAI22X1_30 INVX8_5/A INVX1_47/Y INVX8_2/A INVX2_18/Y gnd OAI22X1_30/Y vdd OAI22X1
XOAI22X1_41 NOR2X1_18/B INVX1_58/Y INVX1_57/Y BUFX4_134/Y gnd NOR2X1_15/B vdd OAI22X1
XFILL_14_6_1 gnd vdd FILL
XOAI22X1_52 OAI22X1_52/A NOR2X1_79/Y NOR2X1_80/Y OAI22X1_52/D gnd OAI22X1_52/Y vdd
+ OAI22X1
XFILL_13_1_0 gnd vdd FILL
XOAI21X1_480 NOR2X1_178/Y MUX2X1_7/A BUFX4_230/Y gnd OAI21X1_480/Y vdd OAI21X1
XOAI22X1_85 MUX2X1_5/B BUFX4_43/Y OAI22X1_85/C OAI22X1_85/D gnd DFFSR_207/D vdd OAI22X1
XOAI22X1_74 OAI22X1_74/A OAI22X1_74/B OAI22X1_74/C OAI22X1_74/D gnd OAI22X1_74/Y vdd
+ OAI22X1
XOAI21X1_491 BUFX4_232/Y OAI21X1_491/B BUFX4_41/Y gnd OAI22X1_98/D vdd OAI21X1
XOAI22X1_96 INVX2_144/Y BUFX4_42/Y OAI22X1_96/C OAI22X1_96/D gnd DFFSR_188/D vdd OAI22X1
XOAI22X1_63 OAI22X1_63/A OAI22X1_63/B OAI22X1_63/C OAI22X1_63/D gnd OAI22X1_63/Y vdd
+ OAI22X1
XFILL_3_3 gnd vdd FILL
XNOR2X1_209 INVX4_12/Y INVX1_152/Y gnd NOR2X1_209/Y vdd NOR2X1
XBUFX4_149 INVX8_23/Y gnd BUFX4_149/Y vdd BUFX4
XBUFX4_138 BUFX4_142/A gnd BUFX4_138/Y vdd BUFX4
XBUFX4_116 BUFX4_117/A gnd BUFX4_116/Y vdd BUFX4
XBUFX4_105 wb_sel_i[0] gnd MUX2X1_41/S vdd BUFX4
XBUFX4_127 DFFSR_245/Q gnd BUFX4_127/Y vdd BUFX4
XFILL_20_4_1 gnd vdd FILL
XFILL_28_5_1 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XINVX2_127 INVX1_56/A gnd MUX2X1_13/A vdd INVX2
XINVX2_105 INVX2_105/A gnd INVX2_105/Y vdd INVX2
XINVX2_138 INVX2_138/A gnd INVX2_138/Y vdd INVX2
XINVX2_149 INVX1_19/A gnd INVX2_149/Y vdd INVX2
XINVX2_116 INVX2_116/A gnd INVX2_116/Y vdd INVX2
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XAOI21X1_186 NOR2X1_209/Y BUFX4_152/Y OAI21X1_555/Y gnd OAI22X1_114/C vdd AOI21X1
XAOI21X1_153 NOR2X1_176/Y BUFX4_152/Y OAI21X1_474/Y gnd OAI22X1_93/C vdd AOI21X1
XAOI21X1_120 INVX2_142/Y OAI21X1_393/B BUFX4_267/Y gnd OAI21X1_393/C vdd AOI21X1
XAOI21X1_142 NOR2X1_170/Y BUFX4_153/Y OAI21X1_434/Y gnd OAI22X1_88/C vdd AOI21X1
XAOI21X1_164 AND2X2_17/Y BUFX4_157/Y OAI21X1_507/Y gnd OAI22X1_102/C vdd AOI21X1
XAOI21X1_175 BUFX4_258/Y OAI21X1_535/Y BUFX4_1/Y gnd AOI22X1_71/D vdd AOI21X1
XAOI21X1_197 INVX2_65/Y OAI21X1_572/B BUFX4_260/Y gnd OAI21X1_572/C vdd AOI21X1
XAOI21X1_131 BUFX4_261/Y OAI21X1_404/Y BUFX4_245/Y gnd AOI22X1_58/D vdd AOI21X1
XOAI22X1_107 INVX2_140/Y BUFX4_166/Y OAI22X1_107/C OAI22X1_107/D gnd DFFSR_172/D vdd
+ OAI22X1
XOAI22X1_118 INVX2_67/Y BUFX4_45/Y OAI22X1_118/C OAI22X1_118/D gnd DFFSR_211/D vdd
+ OAI22X1
XNAND3X1_157 INVX2_66/Y NAND3X1_157/B NAND3X1_157/C gnd NAND3X1_158/C vdd NAND3X1
XNAND3X1_135 INVX2_94/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_137/B vdd NAND3X1
XNAND3X1_113 INVX4_5/Y OAI21X1_217/Y OAI21X1_218/Y gnd NAND3X1_126/B vdd NAND3X1
XNAND3X1_146 INVX1_105/Y BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_148/B vdd NAND3X1
XNAND3X1_102 INVX2_65/Y BUFX4_50/Y BUFX4_136/Y gnd NAND3X1_103/C vdd NAND3X1
XNAND3X1_168 INVX2_107/Y BUFX4_50/Y BUFX4_136/Y gnd NAND3X1_169/C vdd NAND3X1
XNAND3X1_124 INVX2_78/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_125/C vdd NAND3X1
XNAND3X1_179 INVX2_112/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_181/B vdd NAND3X1
XFILL_20_2 gnd vdd FILL
XDFFSR_100 XOR2X1_1/A DFFSR_55/CLK vdd DFFSR_115/S DFFSR_100/D gnd vdd DFFSR
XDFFSR_144 MUX2X1_21/B CLKBUF1_37/Y BUFX4_14/Y vdd DFFSR_144/D gnd vdd DFFSR
XDFFSR_111 NOR3X1_2/A DFFSR_6/CLK vdd DFFSR_113/S DFFSR_111/D gnd vdd DFFSR
XOAI21X1_309 INVX2_72/A NOR2X1_88/B BUFX4_171/Y gnd OAI22X1_69/A vdd OAI21X1
XDFFSR_166 INVX2_122/A CLKBUF1_20/Y BUFX4_12/Y vdd DFFSR_166/D gnd vdd DFFSR
XDFFSR_133 INVX1_103/A CLKBUF1_24/Y BUFX4_13/Y vdd DFFSR_133/D gnd vdd DFFSR
XDFFSR_122 MUX2X1_35/B DFFSR_92/CLK BUFX4_11/Y vdd DFFSR_122/D gnd vdd DFFSR
XBUFX4_7 BUFX4_7/A gnd BUFX4_7/Y vdd BUFX4
XDFFSR_155 INVX2_77/A CLKBUF1_1/Y BUFX4_10/Y vdd DFFSR_155/D gnd vdd DFFSR
XDFFSR_177 INVX2_90/A DFFSR_57/CLK BUFX4_18/Y vdd DFFSR_177/D gnd vdd DFFSR
XDFFSR_188 INVX1_42/A CLKBUF1_41/Y BUFX4_17/Y vdd DFFSR_188/D gnd vdd DFFSR
XDFFSR_199 INVX2_62/A CLKBUF1_6/Y BUFX4_16/Y vdd DFFSR_199/D gnd vdd DFFSR
XFILL_25_3_1 gnd vdd FILL
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XFILL_0_3_1 gnd vdd FILL
XFILL_8_4_1 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_128 BUFX4_28/Y BUFX4_120/Y DFFSR_3/Q gnd BUFX2_5/A vdd OAI21X1
XOAI21X1_117 INVX2_43/Y MUX2X1_35/S OAI21X1_85/C gnd NAND3X1_64/B vdd OAI21X1
XOAI21X1_106 AND2X2_3/Y INVX2_37/Y NAND3X1_58/Y gnd DFFSR_61/D vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd ss_pad_o[1] vdd BUFX2
XOAI21X1_139 BUFX4_27/Y BUFX4_118/Y INVX2_7/A gnd BUFX2_16/A vdd OAI21X1
XNAND2X1_123 AOI21X1_62/B OAI21X1_243/Y gnd OAI21X1_244/B vdd NAND2X1
XNAND2X1_112 INVX4_8/Y OR2X2_6/A gnd AOI22X1_34/A vdd NAND2X1
XNAND2X1_101 MUX2X1_5/Y BUFX4_66/Y gnd AOI21X1_31/B vdd NAND2X1
XNAND2X1_134 NOR2X1_85/A NOR2X1_72/B gnd INVX2_154/A vdd NAND2X1
XNAND2X1_189 NOR2X1_152/Y INVX1_139/A gnd OAI21X1_393/B vdd NAND2X1
XNAND2X1_145 OAI21X1_338/Y OAI21X1_343/Y gnd OAI21X1_344/B vdd NAND2X1
XNAND2X1_167 BUFX4_190/Y wb_dat_i[20] gnd OAI21X1_609/C vdd NAND2X1
XNAND2X1_178 INVX1_141/A INVX8_14/A gnd NAND2X1_178/Y vdd NAND2X1
XNAND2X1_156 INVX1_142/A NOR2X1_71/Y gnd AOI21X1_88/B vdd NAND2X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XOAI21X1_673 NOR2X1_247/Y INVX2_70/Y BUFX4_233/Y gnd OAI21X1_673/Y vdd OAI21X1
XOAI21X1_640 AND2X2_27/Y OAI21X1_640/B OAI21X1_640/C gnd DFFSR_126/D vdd OAI21X1
XAOI21X1_4 INVX1_95/A BUFX4_114/Y AOI21X1_4/C gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_651 INVX1_118/Y BUFX4_111/Y OAI21X1_651/C gnd OAI21X1_651/Y vdd OAI21X1
XOAI21X1_662 BUFX4_163/Y MUX2X1_43/Y OAI21X1_662/C gnd DFFSR_116/D vdd OAI21X1
XOAI21X1_684 BUFX4_121/Y INVX8_20/Y MUX2X1_46/Y gnd OAI21X1_685/C vdd OAI21X1
XXNOR2X1_12 XNOR2X1_9/Y XNOR2X1_12/B gnd XNOR2X1_12/Y vdd XNOR2X1
XOAI21X1_695 INVX1_97/A NOR2X1_251/Y OAI21X1_695/C gnd OAI21X1_696/A vdd OAI21X1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XBUFX2_33 BUFX2_33/A gnd ss_pad_o[30] vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd ss_pad_o[19] vdd BUFX2
XBUFX2_44 DFFSR_73/Q gnd wb_dat_o[8] vdd BUFX2
XBUFX2_11 BUFX2_11/A gnd ss_pad_o[8] vdd BUFX2
XBUFX2_77 INVX1_17/A gnd BUFX2_77/Y vdd BUFX2
XBUFX2_66 DFFSR_95/Q gnd wb_dat_o[30] vdd BUFX2
XBUFX2_55 DFFSR_84/Q gnd wb_dat_o[19] vdd BUFX2
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_23 INVX2_47/Y NOR3X1_1/Y INVX1_74/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_12 INVX1_92/A BUFX4_117/Y OAI22X1_36/Y gnd NAND2X1_46/A vdd AOI21X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_34 AOI21X1_34/A AOI21X1_34/B INVX8_13/Y gnd AOI21X1_34/Y vdd AOI21X1
XAOI21X1_67 AOI21X1_67/A AOI21X1_67/B INVX4_3/Y gnd AOI21X1_68/C vdd AOI21X1
XOAI21X1_7 INVX1_4/Y BUFX4_86/Y OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_56 AOI21X1_56/A AOI21X1_56/B INVX8_13/Y gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_89 BUFX4_265/Y AOI21X1_89/B BUFX4_246/Y gnd AOI22X1_40/D vdd AOI21X1
XAOI21X1_78 INVX2_68/Y AOI21X1_78/B BUFX4_265/Y gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B INVX8_13/Y gnd AOI21X1_45/Y vdd AOI21X1
XFILL_5_2_1 gnd vdd FILL
XOAI22X1_53 OAI22X1_53/A NOR2X1_81/Y NOR2X1_82/Y OAI22X1_53/D gnd OAI22X1_53/Y vdd
+ OAI22X1
XOAI22X1_42 INVX8_5/A INVX1_59/Y INVX8_2/A BUFX4_29/Y gnd OAI22X1_42/Y vdd OAI22X1
XOAI22X1_20 INVX8_1/A INVX2_16/Y INVX2_45/Y INVX8_4/A gnd NOR2X1_8/A vdd OAI22X1
XOAI22X1_31 INVX8_6/A INVX1_49/Y INVX1_48/Y BUFX4_133/Y gnd NOR2X1_12/B vdd OAI22X1
XOAI22X1_64 OAI22X1_64/A OAI22X1_64/B OAI22X1_64/C OAI22X1_64/D gnd OAI22X1_64/Y vdd
+ OAI22X1
XOAI22X1_75 OAI22X1_75/A OAI22X1_75/B OAI22X1_75/C OAI22X1_75/D gnd OAI22X1_75/Y vdd
+ OAI22X1
XFILL_13_1_1 gnd vdd FILL
XOAI21X1_481 MUX2X1_7/A BUFX4_20/Y OAI21X1_641/C gnd OAI21X1_482/B vdd OAI21X1
XOAI21X1_470 BUFX4_232/Y OAI21X1_470/B BUFX4_43/Y gnd OAI22X1_91/D vdd OAI21X1
XOAI22X1_86 INVX2_117/Y BUFX4_42/Y OAI22X1_86/C OAI22X1_86/D gnd DFFSR_206/D vdd OAI22X1
XOAI21X1_492 BUFX4_155/Y OAI21X1_492/B OAI21X1_492/C gnd AOI22X1_68/C vdd OAI21X1
XOAI22X1_97 INVX2_114/Y BUFX4_45/Y OAI22X1_97/C OAI22X1_97/D gnd DFFSR_186/D vdd OAI22X1
XFILL_3_4 gnd vdd FILL
XBUFX4_117 BUFX4_117/A gnd BUFX4_117/Y vdd BUFX4
XBUFX4_128 INVX8_4/Y gnd AND2X2_3/A vdd BUFX4
XBUFX4_139 BUFX4_142/A gnd BUFX4_139/Y vdd BUFX4
XBUFX4_106 wb_sel_i[0] gnd BUFX4_106/Y vdd BUFX4
XFILL_1_1 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XINVX2_128 INVX2_128/A gnd MUX2X1_13/B vdd INVX2
XINVX2_117 INVX2_117/A gnd INVX2_117/Y vdd INVX2
XINVX2_106 INVX2_106/A gnd INVX2_106/Y vdd INVX2
XINVX2_139 INVX2_139/A gnd INVX2_139/Y vdd INVX2
XFILL_18_0_1 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XFILL_21_7_0 gnd vdd FILL
XAOI21X1_110 MUX2X1_9/A OAI21X1_382/B BUFX4_264/Y gnd OAI21X1_382/C vdd AOI21X1
XAOI21X1_121 BUFX4_267/Y OAI21X1_394/Y BUFX4_247/Y gnd AOI22X1_53/D vdd AOI21X1
XAOI21X1_132 INVX2_94/Y OAI21X1_405/B BUFX4_267/Y gnd OAI21X1_405/C vdd AOI21X1
XAOI21X1_165 NOR2X1_190/Y BUFX4_154/Y OAI21X1_510/Y gnd OAI22X1_103/C vdd AOI21X1
XAOI21X1_154 NOR2X1_177/Y BUFX4_154/Y OAI21X1_477/Y gnd OAI22X1_94/C vdd AOI21X1
XAOI21X1_187 INVX2_119/Y OAI21X1_558/B BUFX4_259/Y gnd OAI21X1_558/C vdd AOI21X1
XAOI21X1_176 AND2X2_20/Y BUFX4_157/Y OAI21X1_536/Y gnd OAI22X1_110/C vdd AOI21X1
XAOI21X1_143 INVX2_111/Y OR2X2_11/Y BUFX4_251/Y gnd OAI21X1_438/C vdd AOI21X1
XAOI21X1_198 BUFX4_260/Y OAI21X1_573/Y BUFX4_3/Y gnd AOI22X1_79/D vdd AOI21X1
XOAI22X1_119 INVX2_70/Y BUFX4_42/Y OAI22X1_119/C OAI22X1_119/D gnd DFFSR_195/D vdd
+ OAI22X1
XOAI22X1_108 INVX2_110/Y BUFX4_165/Y OAI22X1_108/C OAI22X1_108/D gnd DFFSR_170/D vdd
+ OAI22X1
XNAND3X1_114 INVX2_73/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_116/B vdd NAND3X1
XNAND3X1_103 BUFX4_206/Y NAND3X1_103/B NAND3X1_103/C gnd AOI21X1_34/B vdd NAND3X1
XNAND3X1_158 INVX4_5/A NAND3X1_158/B NAND3X1_158/C gnd NAND3X1_159/C vdd NAND3X1
XNAND3X1_136 INVX2_95/Y BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_137/C vdd NAND3X1
XNAND3X1_147 INVX2_99/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_148/C vdd NAND3X1
XNAND3X1_169 BUFX4_205/Y NAND3X1_169/B NAND3X1_169/C gnd AOI21X1_45/A vdd NAND3X1
XNAND3X1_125 BUFX4_64/Y NAND3X1_125/B NAND3X1_125/C gnd AOI21X1_40/B vdd NAND3X1
XFILL_12_7_0 gnd vdd FILL
XFILL_20_3 gnd vdd FILL
XDFFSR_101 XOR2X1_1/B DFFSR_41/CLK vdd DFFSR_99/R DFFSR_101/D gnd vdd DFFSR
XDFFSR_189 INVX2_81/A CLKBUF1_37/Y BUFX4_15/Y vdd DFFSR_189/D gnd vdd DFFSR
XDFFSR_112 NOR2X1_22/B DFFSR_7/CLK vdd DFFSR_113/S DFFSR_112/D gnd vdd DFFSR
XBUFX4_8 BUFX4_9/A gnd BUFX4_8/Y vdd BUFX4
XDFFSR_156 INVX1_43/A CLKBUF1_49/Y BUFX4_18/Y vdd DFFSR_156/D gnd vdd DFFSR
XDFFSR_178 INVX2_104/A CLKBUF1_24/Y BUFX4_13/Y vdd DFFSR_178/D gnd vdd DFFSR
XDFFSR_167 INVX2_61/A CLKBUF1_15/Y BUFX4_13/Y vdd DFFSR_167/D gnd vdd DFFSR
XDFFSR_134 INVX1_114/A CLKBUF1_6/A BUFX4_13/Y vdd DFFSR_134/D gnd vdd DFFSR
XDFFSR_123 INVX1_99/A DFFSR_3/CLK BUFX4_11/Y vdd DFFSR_123/D gnd vdd DFFSR
XDFFSR_145 MUX2X1_19/B DFFSR_85/CLK BUFX4_11/Y vdd DFFSR_145/D gnd vdd DFFSR
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XOAI21X1_129 BUFX4_27/Y BUFX4_118/Y DFFSR_4/Q gnd BUFX2_6/A vdd OAI21X1
XOAI21X1_107 INVX2_38/Y BUFX4_24/Y OAI21X1_47/C gnd NAND3X1_59/B vdd OAI21X1
XOAI21X1_118 AND2X2_3/Y INVX2_43/Y NAND3X1_64/Y gnd DFFSR_51/D vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd ss_pad_o[2] vdd BUFX2
XNAND2X1_124 OAI21X1_241/C AOI21X1_69/B gnd INVX1_129/A vdd NAND2X1
XNAND2X1_135 AOI22X1_34/B AOI22X1_34/A gnd OAI21X1_256/C vdd NAND2X1
XNAND2X1_113 OR2X2_5/A OR2X2_5/B gnd OAI21X1_235/A vdd NAND2X1
XNAND2X1_102 BUFX4_183/Y OR2X2_6/A gnd BUFX4_76/A vdd NAND2X1
XNAND2X1_179 NOR2X1_147/Y INVX1_139/A gnd OAI21X1_382/B vdd NAND2X1
XNAND2X1_146 OAI21X1_323/Y OAI21X1_344/Y gnd OAI21X1_345/B vdd NAND2X1
XNAND2X1_168 NOR2X1_156/Y NOR2X1_71/Y gnd OAI21X1_370/B vdd NAND2X1
XNAND2X1_157 BUFX4_91/Y wb_dat_i[26] gnd OAI21X1_520/C vdd NAND2X1
XFILL_26_6_0 gnd vdd FILL
XNOR2X1_190 INVX4_11/Y INVX1_150/Y gnd NOR2X1_190/Y vdd NOR2X1
XFILL_1_6_0 gnd vdd FILL
XOAI21X1_641 INVX1_100/Y BUFX4_26/Y OAI21X1_641/C gnd OAI21X1_641/Y vdd OAI21X1
XOAI21X1_630 MUX2X1_12/A BUFX4_22/Y OAI21X1_630/C gnd OAI21X1_630/Y vdd OAI21X1
XOAI21X1_674 INVX2_70/Y BUFX4_22/Y OAI21X1_694/C gnd OAI21X1_675/B vdd OAI21X1
XOAI21X1_663 BUFX4_55/Y BUFX4_125/Y NOR2X1_75/Y gnd NOR2X1_247/B vdd OAI21X1
XOAI21X1_696 OAI21X1_696/A BUFX4_4/Y OAI21X1_696/C gnd DFFSR_131/D vdd OAI21X1
XOAI21X1_652 INVX1_118/A NOR2X1_239/Y OAI21X1_652/C gnd OAI21X1_653/A vdd OAI21X1
XAOI21X1_5 INVX1_118/A BUFX4_113/Y AOI21X1_5/C gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_685 BUFX4_163/Y MUX2X1_45/Y OAI21X1_685/C gnd DFFSR_147/D vdd OAI21X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XXNOR2X1_13 XNOR2X1_13/A OR2X2_8/Y gnd XNOR2X1_13/Y vdd XNOR2X1
XFILL_9_7_0 gnd vdd FILL
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XBUFX2_78 INVX4_8/A gnd BUFX2_78/Y vdd BUFX2
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XBUFX2_45 DFFSR_74/Q gnd wb_dat_o[9] vdd BUFX2
XINVX1_92 INVX1_92/A gnd MUX2X1_3/A vdd INVX1
XFILL_17_6_0 gnd vdd FILL
XBUFX2_34 BUFX2_34/A gnd ss_pad_o[31] vdd BUFX2
XBUFX2_56 DFFSR_85/Q gnd wb_dat_o[20] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd ss_pad_o[20] vdd BUFX2
XBUFX2_67 DFFSR_96/Q gnd wb_dat_o[31] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd ss_pad_o[9] vdd BUFX2
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_68 OR2X2_8/Y AOI21X1_68/B AOI21X1_68/C gnd XNOR2X1_12/B vdd AOI21X1
XAOI21X1_24 INVX1_75/A NOR3X1_1/Y INVX1_76/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_13 MUX2X1_33/B BUFX4_117/Y OAI22X1_39/Y gnd NAND2X1_47/A vdd AOI21X1
XAOI21X1_57 AOI21X1_57/A AOI21X1_57/B BUFX4_81/Y gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B BUFX4_81/Y gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_35 AOI21X1_35/A AOI21X1_35/B BUFX4_205/Y gnd AOI21X1_35/Y vdd AOI21X1
XOAI21X1_8 OAI21X1_8/A INVX1_4/Y OAI21X1_8/C gnd DFFSR_28/D vdd OAI21X1
XAOI21X1_79 BUFX4_265/Y AOI21X1_79/B BUFX4_246/Y gnd AOI22X1_35/D vdd AOI21X1
XOAI22X1_87 MUX2X1_7/B BUFX4_44/Y OAI22X1_87/C OAI22X1_87/D gnd DFFSR_205/D vdd OAI22X1
XOAI22X1_54 OAI22X1_54/A NOR2X1_83/Y NOR2X1_84/Y OAI22X1_54/D gnd OAI22X1_54/Y vdd
+ OAI22X1
XOAI22X1_32 BUFX4_193/Y INVX2_4/Y INVX2_33/Y BUFX4_220/Y gnd NOR2X1_12/A vdd OAI22X1
XOAI22X1_98 INVX2_102/Y BUFX4_41/Y OAI22X1_98/C OAI22X1_98/D gnd DFFSR_185/D vdd OAI22X1
XOAI22X1_65 OAI22X1_65/A OAI22X1_65/B OAI22X1_65/C OAI22X1_65/D gnd OAI22X1_65/Y vdd
+ OAI22X1
XOAI22X1_10 INVX8_6/A INVX1_28/Y INVX1_27/Y BUFX4_133/Y gnd NOR2X1_5/B vdd OAI22X1
XOAI22X1_76 OAI22X1_76/A OAI22X1_76/B OAI22X1_76/C OAI22X1_76/D gnd OAI22X1_76/Y vdd
+ OAI22X1
XOAI22X1_43 OAI22X1_8/D INVX2_37/Y OAI22X1_7/A INVX1_60/Y gnd OAI22X1_43/Y vdd OAI22X1
XOAI22X1_21 INVX8_5/A INVX1_38/Y INVX8_2/A INVX2_29/Y gnd AOI21X1_7/C vdd OAI22X1
XOAI21X1_482 BUFX4_230/Y OAI21X1_482/B BUFX4_44/Y gnd OAI22X1_95/D vdd OAI21X1
XOAI21X1_471 NOR2X1_175/Y MUX2X1_14/A BUFX4_230/Y gnd OAI21X1_471/Y vdd OAI21X1
XOAI21X1_460 BUFX4_146/Y OAI21X1_460/B BUFX4_249/Y gnd AOI22X1_65/D vdd OAI21X1
XOAI21X1_493 INVX2_135/Y MUX2X1_41/S OAI21X1_651/C gnd OAI21X1_494/B vdd OAI21X1
XFILL_23_4_0 gnd vdd FILL
XBUFX4_118 DFFSR_245/Q gnd BUFX4_118/Y vdd BUFX4
XFILL_6_5_0 gnd vdd FILL
XBUFX4_107 wb_sel_i[0] gnd MUX2X1_43/S vdd BUFX4
XBUFX4_129 INVX8_4/Y gnd BUFX4_129/Y vdd BUFX4
XFILL_14_4_0 gnd vdd FILL
XOAI21X1_290 NOR2X1_82/B MUX2X1_21/B BUFX4_33/Y gnd OAI22X1_62/D vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XINVX2_129 INVX1_54/A gnd MUX2X1_14/A vdd INVX2
XDFFSR_90 DFFSR_90/Q CLKBUF1_3/A DFFSR_2/R vdd DFFSR_90/D gnd vdd DFFSR
XINVX2_107 INVX1_60/A gnd INVX2_107/Y vdd INVX2
XINVX2_118 INVX1_50/A gnd INVX2_118/Y vdd INVX2
XFILL_30_7_1 gnd vdd FILL
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XAOI21X1_155 NOR2X1_178/Y BUFX4_152/Y OAI21X1_480/Y gnd OAI22X1_95/C vdd AOI21X1
XAOI21X1_166 NOR2X1_192/Y BUFX4_152/Y OAI21X1_513/Y gnd OAI22X1_104/C vdd AOI21X1
XFILL_21_7_1 gnd vdd FILL
XAOI21X1_111 BUFX4_263/Y OAI21X1_383/Y BUFX4_243/Y gnd AOI22X1_49/D vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XAOI21X1_133 BUFX4_267/Y OAI21X1_406/Y BUFX4_247/Y gnd AOI22X1_59/D vdd AOI21X1
XAOI21X1_122 INVX2_112/Y OAI21X1_395/B BUFX4_268/Y gnd OAI21X1_395/C vdd AOI21X1
XAOI21X1_100 INVX2_60/Y OAI21X1_370/B BUFX4_262/Y gnd OAI21X1_370/C vdd AOI21X1
XAOI21X1_144 NOR2X1_171/Y BUFX4_159/Y OAI21X1_442/Y gnd OAI22X1_89/C vdd AOI21X1
XAOI21X1_188 BUFX4_259/Y OAI21X1_559/Y BUFX4_4/Y gnd AOI22X1_75/D vdd AOI21X1
XAOI21X1_177 INVX2_122/Y OAI21X1_539/B BUFX4_258/Y gnd OAI21X1_539/C vdd AOI21X1
XAOI21X1_199 INVX2_125/Y OAI21X1_574/B BUFX4_260/Y gnd OAI21X1_574/C vdd AOI21X1
XFILL_28_3_0 gnd vdd FILL
XOAI22X1_109 INVX2_98/Y BUFX4_161/Y OAI22X1_109/C OAI22X1_109/D gnd DFFSR_169/D vdd
+ OAI22X1
XNAND3X1_104 NOR3X1_4/B OAI21X1_214/Y OAI21X1_216/Y gnd NAND3X1_127/B vdd NAND3X1
XNAND3X1_126 INVX2_66/Y NAND3X1_126/B OAI21X1_219/Y gnd NAND3X1_127/C vdd NAND3X1
XNAND3X1_137 BUFX4_207/Y NAND3X1_137/B NAND3X1_137/C gnd NAND3X1_141/B vdd NAND3X1
XFILL_3_3_0 gnd vdd FILL
XNAND3X1_115 INVX2_74/Y BUFX4_51/Y BUFX4_141/Y gnd NAND3X1_116/C vdd NAND3X1
XNAND3X1_148 BUFX4_64/Y NAND3X1_148/B NAND3X1_148/C gnd NAND3X1_149/C vdd NAND3X1
XNAND3X1_159 INVX1_86/A OAI21X1_223/Y NAND3X1_159/C gnd NAND3X1_160/B vdd NAND3X1
XFILL_11_2_0 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFSR_157 INVX2_79/A DFFSR_37/CLK BUFX4_15/Y vdd DFFSR_157/D gnd vdd DFFSR
XDFFSR_113 NOR3X1_3/A DFFSR_8/CLK vdd DFFSR_113/S DFFSR_113/D gnd vdd DFFSR
XDFFSR_102 INVX1_68/A DFFSR_57/CLK vdd DFFSR_108/S DFFSR_102/D gnd vdd DFFSR
XDFFSR_124 INVX1_121/A CLKBUF1_5/Y BUFX4_18/Y vdd DFFSR_124/D gnd vdd DFFSR
XDFFSR_168 INVX2_137/A CLKBUF1_10/Y BUFX4_12/Y vdd DFFSR_168/D gnd vdd DFFSR
XDFFSR_146 MUX2X1_17/B DFFSR_86/CLK BUFX4_13/Y vdd DFFSR_146/D gnd vdd DFFSR
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XDFFSR_135 INVX1_94/A CLKBUF1_6/A BUFX4_10/Y vdd DFFSR_135/D gnd vdd DFFSR
XDFFSR_179 INVX2_69/A CLKBUF1_6/A BUFX4_10/Y vdd DFFSR_179/D gnd vdd DFFSR
XINVX4_9 INVX4_9/A gnd INVX4_9/Y vdd INVX4
XNAND3X1_90 INVX1_72/Y AND2X2_4/Y AND2X2_5/Y gnd NOR3X1_3/C vdd NAND3X1
XNOR2X1_90 INVX2_79/A NOR2X1_99/B gnd NOR2X1_90/Y vdd NOR2X1
XOAI21X1_119 INVX2_44/Y MUX2X1_37/S OAI21X1_87/C gnd NAND3X1_65/B vdd OAI21X1
XOAI21X1_108 AND2X2_3/Y INVX2_38/Y NAND3X1_59/Y gnd DFFSR_62/D vdd OAI21X1
XNAND2X1_114 INVX4_8/A OR2X2_7/B gnd OAI21X1_251/C vdd NAND2X1
XNAND2X1_125 INVX4_8/Y AND2X2_10/Y gnd OAI21X1_247/C vdd NAND2X1
XNAND2X1_103 INVX1_100/Y MUX2X1_6/S gnd OAI21X1_220/C vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd ss_pad_o[3] vdd BUFX2
XNAND2X1_158 NOR2X1_151/Y NOR2X1_71/Y gnd AOI21X1_90/B vdd NAND2X1
XNAND2X1_136 OAI21X1_263/Y OAI21X1_268/Y gnd OAI21X1_279/A vdd NAND2X1
XNAND2X1_169 BUFX4_185/Y wb_dat_i[19] gnd OAI21X1_613/C vdd NAND2X1
XNAND2X1_1 wb_dat_i[24] BUFX4_86/Y gnd OAI21X1_1/C vdd NAND2X1
XNAND2X1_147 wb_dat_i[31] BUFX4_88/Y gnd OAI21X1_672/C vdd NAND2X1
XFILL_26_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XNOR2X1_191 INVX8_18/A NOR2X1_191/B gnd INVX1_151/A vdd NOR2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XFILL_1_6_1 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_180 INVX8_19/Y OR2X2_11/A gnd NOR2X1_180/Y vdd NOR2X1
XOAI21X1_642 AND2X2_28/B INVX1_100/A MUX2X1_26/S gnd OAI21X1_643/B vdd OAI21X1
XOAI21X1_631 AND2X2_25/B INVX1_101/A BUFX4_162/Y gnd OAI21X1_632/B vdd OAI21X1
XAOI21X1_6 MUX2X1_37/B BUFX4_115/Y AOI21X1_6/C gnd AOI21X1_6/Y vdd AOI21X1
XOAI21X1_675 BUFX4_233/Y OAI21X1_675/B BUFX4_42/Y gnd OAI22X1_119/D vdd OAI21X1
XOAI21X1_686 BUFX4_153/Y OAI21X1_686/B OAI21X1_686/C gnd AOI22X1_86/C vdd OAI21X1
XOAI21X1_664 NOR2X1_244/Y INVX2_67/Y BUFX4_229/Y gnd OAI21X1_664/Y vdd OAI21X1
XOAI21X1_697 INVX1_98/Y BUFX4_190/Y OAI21X1_697/C gnd OAI21X1_697/Y vdd OAI21X1
XOAI21X1_620 AND2X2_24/Y OAI21X1_620/B OAI21X1_620/C gnd DFFSR_134/D vdd OAI21X1
XOAI21X1_653 OAI21X1_653/A BUFX4_2/Y OAI21X1_653/C gnd DFFSR_120/D vdd OAI21X1
XXNOR2X1_14 OR2X2_5/A INVX4_9/A gnd XNOR2X1_14/Y vdd XNOR2X1
XFILL_8_2_0 gnd vdd FILL
XFILL_9_7_1 gnd vdd FILL
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XINVX1_82 BUFX2_1/A gnd INVX1_82/Y vdd INVX1
XBUFX2_79 MUX2X1_1/S gnd BUFX2_79/Y vdd BUFX2
XINVX1_71 INVX2_31/A gnd INVX1_71/Y vdd INVX1
XBUFX2_35 DFFSR_64/Q gnd wb_ack_o vdd BUFX2
XINVX1_93 INVX1_93/A gnd MUX2X1_3/B vdd INVX1
XBUFX2_13 BUFX2_13/A gnd ss_pad_o[10] vdd BUFX2
XFILL_17_6_1 gnd vdd FILL
XFILL_16_1_0 gnd vdd FILL
XBUFX2_46 DFFSR_75/Q gnd wb_dat_o[10] vdd BUFX2
XBUFX2_68 gnd gnd wb_err_o vdd BUFX2
XBUFX2_24 BUFX2_24/A gnd ss_pad_o[21] vdd BUFX2
XBUFX2_57 DFFSR_86/Q gnd wb_dat_o[21] vdd BUFX2
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_69 INVX2_151/Y AOI21X1_69/B NOR3X1_7/B gnd AOI21X1_69/Y vdd AOI21X1
XAOI21X1_25 INVX1_78/Y NOR3X1_1/Y INVX1_77/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_14 INVX1_101/A BUFX4_115/Y OAI22X1_42/Y gnd NAND2X1_48/A vdd AOI21X1
XAOI21X1_36 AOI21X1_36/A AOI21X1_36/B BUFX4_65/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_58 AOI21X1_58/A AOI21X1_58/B INVX8_13/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_47 AOI21X1_47/A AOI21X1_47/B INVX8_13/Y gnd AOI21X1_47/Y vdd AOI21X1
XOAI21X1_9 INVX1_5/Y BUFX4_88/Y OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_88 INVX2_141/Y BUFX4_41/Y OAI22X1_88/C OAI22X1_88/D gnd DFFSR_204/D vdd OAI22X1
XOAI22X1_11 OAI22X1_5/A INVX2_13/Y INVX2_42/Y OAI22X1_5/D gnd NOR2X1_5/A vdd OAI22X1
XOAI22X1_66 OAI22X1_66/A OAI22X1_66/B OAI22X1_66/C OAI22X1_66/D gnd OAI22X1_66/Y vdd
+ OAI22X1
XOAI22X1_33 INVX8_5/A INVX1_50/Y INVX8_2/A INVX2_20/Y gnd OAI22X1_33/Y vdd OAI22X1
XOAI22X1_55 OAI22X1_55/A NOR2X1_86/Y NOR2X1_87/Y OAI22X1_55/D gnd OAI22X1_55/Y vdd
+ OAI22X1
XOAI22X1_77 OAI22X1_77/A OAI22X1_77/B OAI22X1_77/C OAI22X1_77/D gnd OAI22X1_77/Y vdd
+ OAI22X1
XOAI21X1_450 NOR2X1_172/Y INVX2_62/Y BUFX4_229/Y gnd OAI21X1_450/Y vdd OAI21X1
XOAI22X1_44 OAI22X1_8/A INVX2_8/Y BUFX4_133/Y INVX1_61/Y gnd OAI22X1_44/Y vdd OAI22X1
XOAI22X1_22 INVX8_6/A INVX1_40/Y INVX1_39/Y BUFX4_133/Y gnd NOR2X1_9/B vdd OAI22X1
XOAI22X1_99 INVX2_63/Y BUFX4_45/Y OAI22X1_99/C OAI22X1_99/D gnd DFFSR_183/D vdd OAI22X1
XOAI21X1_472 MUX2X1_14/A BUFX4_25/Y OAI21X1_553/C gnd OAI21X1_473/B vdd OAI21X1
XOAI21X1_483 NOR2X1_179/Y INVX2_144/Y BUFX4_233/Y gnd OAI21X1_483/Y vdd OAI21X1
XOAI21X1_494 BUFX4_144/Y OAI21X1_494/B BUFX4_248/Y gnd AOI22X1_68/D vdd OAI21X1
XOAI21X1_461 BUFX4_54/Y BUFX4_126/Y NOR2X1_160/Y gnd INVX1_148/A vdd OAI21X1
XFILL_23_4_1 gnd vdd FILL
XBUFX4_119 DFFSR_245/Q gnd INVX4_10/A vdd BUFX4
XFILL_5_0_0 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XBUFX4_108 wb_sel_i[0] gnd BUFX4_108/Y vdd BUFX4
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_280 INVX4_9/Y INVX4_8/A OAI21X1_280/C gnd OAI21X1_281/C vdd OAI21X1
XOAI21X1_291 OAI22X1_61/Y OAI22X1_62/Y NOR2X1_72/Y gnd OAI21X1_291/Y vdd OAI21X1
XFILL_1_3 gnd vdd FILL
XFILL_29_1 gnd vdd FILL
XINVX2_119 INVX1_49/A gnd INVX2_119/Y vdd INVX2
XINVX2_108 INVX1_61/A gnd INVX2_108/Y vdd INVX2
XDFFSR_80 DFFSR_80/Q CLKBUF1_3/Y DFFSR_80/R vdd DFFSR_80/D gnd vdd DFFSR
XDFFSR_91 DFFSR_91/Q DFFSR_91/CLK DFFSR_9/R vdd DFFSR_91/D gnd vdd DFFSR
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_130 BUFX4_78/Y gnd NOR2X1_71/B vdd INVX1
XINVX1_141 INVX1_141/A gnd INVX1_141/Y vdd INVX1
XAOI21X1_189 NOR2X1_210/Y BUFX4_152/Y OAI21X1_560/Y gnd OAI22X1_115/C vdd AOI21X1
XAOI21X1_167 NOR2X1_194/Y BUFX4_152/Y OAI21X1_516/Y gnd OAI22X1_105/C vdd AOI21X1
XAOI21X1_112 MUX2X1_13/A OAI21X1_384/B BUFX4_264/Y gnd OAI21X1_384/C vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_156 NOR2X1_179/Y BUFX4_156/Y OAI21X1_483/Y gnd OAI22X1_96/C vdd AOI21X1
XAOI21X1_123 BUFX4_268/Y OAI21X1_396/Y BUFX4_247/Y gnd AOI22X1_54/D vdd AOI21X1
XAOI21X1_178 BUFX4_258/Y OAI21X1_540/Y BUFX4_1/Y gnd AOI22X1_72/D vdd AOI21X1
XAOI21X1_145 INVX2_138/Y OAI21X1_446/B BUFX4_255/Y gnd OAI21X1_446/C vdd AOI21X1
XAOI21X1_101 BUFX4_262/Y OAI21X1_371/Y BUFX4_248/Y gnd AOI22X1_46/D vdd AOI21X1
XAOI21X1_134 INVX2_148/Y OAI21X1_407/B BUFX4_261/Y gnd OAI21X1_407/C vdd AOI21X1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XNAND3X1_127 INVX1_86/Y NAND3X1_127/B NAND3X1_127/C gnd NAND3X1_160/C vdd NAND3X1
XNAND3X1_138 INVX1_104/Y BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_140/B vdd NAND3X1
XNAND3X1_116 BUFX4_204/Y NAND3X1_116/B NAND3X1_116/C gnd AOI21X1_39/A vdd NAND3X1
XNAND3X1_149 INVX8_13/Y NAND3X1_149/B NAND3X1_149/C gnd NAND3X1_157/B vdd NAND3X1
XNAND3X1_105 INVX1_96/Y BUFX4_50/Y BUFX4_137/Y gnd AOI21X1_35/A vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFSR_114 NOR2X1_23/B DFFSR_99/CLK vdd DFFSR_115/S DFFSR_114/D gnd vdd DFFSR
XDFFSR_103 NOR2X1_28/A DFFSR_58/CLK vdd DFFSR_108/S DFFSR_103/D gnd vdd DFFSR
XDFFSR_125 INVX1_100/A CLKBUF1_2/Y BUFX4_14/Y vdd DFFSR_125/D gnd vdd DFFSR
XDFFSR_136 INVX1_119/A CLKBUF1_19/Y BUFX4_16/Y vdd DFFSR_136/D gnd vdd DFFSR
XDFFSR_169 INVX2_98/A CLKBUF1_6/Y BUFX4_13/Y vdd DFFSR_169/D gnd vdd DFFSR
XDFFSR_147 INVX1_96/A CLKBUF1_25/Y BUFX4_11/Y vdd DFFSR_147/D gnd vdd DFFSR
XDFFSR_158 INVX1_49/A DFFSR_83/CLK BUFX4_11/Y vdd DFFSR_158/D gnd vdd DFFSR
XNAND3X1_91 XOR2X1_4/B XOR2X1_5/B XOR2X1_4/A gnd NAND3X1_91/Y vdd NAND3X1
XNAND3X1_80 NAND3X1_80/A NAND3X1_80/B NAND3X1_80/C gnd DFFSR_89/D vdd NAND3X1
XNOR2X1_91 INVX2_80/A NOR2X1_99/B gnd NOR2X1_91/Y vdd NOR2X1
XNOR2X1_80 INVX2_91/A NOR2X1_89/B gnd NOR2X1_80/Y vdd NOR2X1
XOAI21X1_109 INVX2_39/Y MUX2X1_41/S OAI21X1_77/C gnd NAND3X1_60/B vdd OAI21X1
XFILL_11_1 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd ss_pad_o[4] vdd BUFX2
XNAND2X1_126 OAI21X1_236/Y XNOR2X1_9/Y gnd OAI21X1_249/C vdd NAND2X1
XNAND2X1_115 OR2X2_5/B INVX4_8/Y gnd AOI21X1_63/A vdd NAND2X1
XNAND2X1_159 BUFX4_86/Y wb_dat_i[25] gnd OAI21X1_522/C vdd NAND2X1
XNAND2X1_104 MUX2X1_9/Y NOR2X1_66/B gnd AOI21X1_42/A vdd NAND2X1
XNAND2X1_137 NOR2X1_85/A NOR2X1_85/B gnd INVX2_155/A vdd NAND2X1
XNAND2X1_148 INVX1_140/A NOR2X1_71/Y gnd AOI21X1_80/B vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XNAND2X1_2 BUFX4_88/Y wb_dat_i[25] gnd OAI21X1_3/C vdd NAND2X1
XNOR2X1_192 INVX4_11/Y INVX1_151/Y gnd NOR2X1_192/Y vdd NOR2X1
XOAI21X1_632 AND2X2_25/Y OAI21X1_632/B OAI21X1_632/C gnd DFFSR_129/D vdd OAI21X1
XNOR2X1_170 OR2X2_13/B NOR2X1_198/B gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_181 INVX8_19/Y NOR2X1_201/B gnd NOR2X1_181/Y vdd NOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XOAI21X1_621 INVX1_103/Y NAND2X1_9/B OAI21X1_621/C gnd OAI21X1_621/Y vdd OAI21X1
XFILL_0_1_1 gnd vdd FILL
XOAI21X1_610 BUFX4_127/Y INVX8_22/Y INVX1_155/Y gnd NOR2X1_239/B vdd OAI21X1
XOAI21X1_643 AND2X2_28/Y OAI21X1_643/B OAI21X1_643/C gnd DFFSR_125/D vdd OAI21X1
XOAI21X1_687 INVX2_71/Y BUFX4_23/Y OAI21X1_694/C gnd OAI21X1_687/Y vdd OAI21X1
XOAI21X1_665 INVX2_67/Y BUFX4_90/Y OAI21X1_672/C gnd OAI21X1_666/B vdd OAI21X1
XOAI21X1_698 BUFX4_127/Y INVX8_22/Y NOR2X1_250/Y gnd NOR2X1_253/B vdd OAI21X1
XAOI21X1_7 MUX2X1_35/B BUFX4_113/Y AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_676 BUFX4_53/Y BUFX4_126/Y NOR2X1_245/Y gnd OR2X2_13/A vdd OAI21X1
XOAI21X1_654 BUFX4_121/Y INVX8_20/Y MUX2X1_40/Y gnd OAI21X1_655/C vdd OAI21X1
XINVX1_72 NOR3X1_1/B gnd INVX1_72/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XFILL_8_2_1 gnd vdd FILL
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XBUFX2_47 DFFSR_76/Q gnd wb_dat_o[11] vdd BUFX2
XBUFX2_36 DFFSR_65/Q gnd wb_dat_o[0] vdd BUFX2
XBUFX2_69 INVX1_64/A gnd wb_int_o vdd BUFX2
XFILL_16_1_1 gnd vdd FILL
XBUFX2_58 DFFSR_87/Q gnd wb_dat_o[22] vdd BUFX2
XBUFX2_14 BUFX2_14/A gnd ss_pad_o[11] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd ss_pad_o[22] vdd BUFX2
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_26 INVX1_80/A NOR2X1_46/A NOR2X1_46/B gnd AOI21X1_27/B vdd AOI21X1
XAOI21X1_59 AOI21X1_59/A AOI21X1_59/B INVX2_66/Y gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_37 AOI21X1_37/A AOI21X1_37/B BUFX4_207/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B INVX8_13/A gnd AOI21X1_48/Y vdd AOI21X1
XAOI21X1_15 INVX2_106/A BUFX4_70/Y OAI22X1_43/Y gnd NAND2X1_49/A vdd AOI21X1
XOAI22X1_34 NOR2X1_18/B INVX1_52/Y INVX1_51/Y BUFX4_134/Y gnd NOR2X1_13/B vdd OAI22X1
XOAI22X1_12 INVX8_5/A INVX1_29/Y INVX8_2/A INVX2_26/Y gnd AOI21X1_4/C vdd OAI22X1
XOAI22X1_23 INVX8_1/A INVX2_17/Y INVX2_46/Y INVX8_4/A gnd NOR2X1_9/A vdd OAI22X1
XOAI21X1_473 BUFX4_230/Y OAI21X1_473/B BUFX4_44/Y gnd OAI22X1_92/D vdd OAI21X1
XOAI21X1_484 INVX2_144/Y BUFX4_21/Y OAI21X1_644/C gnd OAI21X1_485/B vdd OAI21X1
XOAI22X1_56 OAI22X1_56/A NOR2X1_88/Y NOR2X1_89/Y OAI22X1_56/D gnd OAI22X1_56/Y vdd
+ OAI22X1
XOAI22X1_45 OAI22X1_8/D INVX2_38/Y OAI22X1_4/A INVX1_62/Y gnd OAI22X1_45/Y vdd OAI22X1
XOAI21X1_440 BUFX4_145/Y OAI21X1_440/B BUFX4_244/Y gnd AOI22X1_62/D vdd OAI21X1
XOAI21X1_462 BUFX4_158/Y OAI21X1_462/B OAI21X1_462/C gnd AOI22X1_66/C vdd OAI21X1
XOAI22X1_67 OAI22X1_67/A OAI22X1_67/B OAI22X1_67/C OAI22X1_67/D gnd OAI22X1_67/Y vdd
+ OAI22X1
XOAI22X1_89 INVX2_99/Y INVX8_16/A OAI22X1_89/C OAI22X1_89/D gnd DFFSR_201/D vdd OAI22X1
XOAI21X1_451 INVX2_62/Y BUFX4_189/Y OAI21X1_613/C gnd OAI21X1_452/B vdd OAI21X1
XOAI22X1_78 OAI22X1_78/A OAI22X1_78/B OAI22X1_78/C OAI22X1_78/D gnd OAI22X1_78/Y vdd
+ OAI22X1
XOAI21X1_495 NOR2X1_182/Y INVX2_63/Y BUFX4_234/Y gnd OAI21X1_495/Y vdd OAI21X1
XFILL_5_0_1 gnd vdd FILL
XBUFX4_109 wb_sel_i[0] gnd MUX2X1_35/S vdd BUFX4
XOAI21X1_281 INVX1_136/Y OR2X2_1/B OAI21X1_281/C gnd OR2X2_10/A vdd OAI21X1
XOAI21X1_292 INVX1_32/A BUFX4_222/Y BUFX4_169/Y gnd OAI22X1_63/A vdd OAI21X1
XOAI21X1_270 INVX2_97/A NOR2X1_89/B BUFX4_78/Y gnd OAI22X1_55/D vdd OAI21X1
XFILL_29_2 gnd vdd FILL
XFILL_24_7_0 gnd vdd FILL
XINVX2_109 INVX2_109/A gnd INVX2_109/Y vdd INVX2
XDFFSR_70 DFFSR_70/Q DFFSR_70/CLK DFFSR_93/R vdd DFFSR_70/D gnd vdd DFFSR
XDFFSR_81 DFFSR_81/Q DFFSR_96/CLK DFFSR_96/R vdd DFFSR_81/D gnd vdd DFFSR
XDFFSR_92 DFFSR_92/Q DFFSR_92/CLK DFFSR_3/R vdd DFFSR_92/D gnd vdd DFFSR
XFILL_15_7_0 gnd vdd FILL
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_120 MUX2X1_27/B gnd MUX2X1_28/B vdd INVX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XAOI21X1_113 BUFX4_264/Y OAI21X1_385/Y BUFX4_250/Y gnd AOI22X1_50/D vdd AOI21X1
XAOI21X1_124 INVX2_100/Y OAI21X1_397/B BUFX4_267/Y gnd OAI21X1_397/C vdd AOI21X1
XAOI21X1_179 NOR2X1_204/Y BUFX4_157/Y OAI21X1_542/Y gnd OAI22X1_111/C vdd AOI21X1
XAOI21X1_102 INVX2_121/Y INVX1_137/A BUFX4_266/Y gnd AOI21X1_103/A vdd AOI21X1
XAOI21X1_135 BUFX4_261/Y OAI21X1_408/Y BUFX4_245/Y gnd AOI22X1_60/D vdd AOI21X1
XAOI21X1_146 NOR2X1_172/Y BUFX4_159/Y OAI21X1_450/Y gnd OAI22X1_90/C vdd AOI21X1
XAOI21X1_157 NOR2X1_180/Y BUFX4_160/Y OAI21X1_486/Y gnd OAI22X1_97/C vdd AOI21X1
XAOI21X1_168 INVX2_116/Y OAI21X1_519/B BUFX4_257/Y gnd OAI21X1_519/C vdd AOI21X1
XNAND3X1_139 INVX2_96/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_140/C vdd NAND3X1
XNAND3X1_128 INVX1_103/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_130/B vdd NAND3X1
XNAND3X1_117 INVX1_98/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_119/B vdd NAND3X1
XNAND3X1_106 INVX2_67/Y BUFX4_76/Y BUFX4_57/Y gnd AOI21X1_35/B vdd NAND3X1
XFILL_30_5_0 gnd vdd FILL
XDFFSR_104 INVX1_70/A CLKBUF1_5/A vdd DFFSR_115/S DFFSR_104/D gnd vdd DFFSR
XDFFSR_115 INVX1_79/A DFFSR_55/CLK vdd DFFSR_115/S DFFSR_115/D gnd vdd DFFSR
XDFFSR_126 INVX1_113/A CLKBUF1_49/Y BUFX4_18/Y vdd DFFSR_126/D gnd vdd DFFSR
XDFFSR_137 INVX1_105/A CLKBUF1_15/Y BUFX4_13/Y vdd DFFSR_137/D gnd vdd DFFSR
XDFFSR_148 INVX1_19/A CLKBUF1_24/Y BUFX4_16/Y vdd DFFSR_148/D gnd vdd DFFSR
XDFFSR_159 INVX2_53/A CLKBUF1_37/Y BUFX4_14/Y vdd DFFSR_159/D gnd vdd DFFSR
XBUFX4_270 DFFSR_44/Q gnd OR2X2_9/B vdd BUFX4
XFILL_21_5_0 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_4_6_0 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XNAND3X1_81 NAND3X1_81/A NAND3X1_81/B NAND3X1_81/C gnd DFFSR_90/D vdd NAND3X1
XNAND3X1_70 INVX4_1/Y INVX2_1/Y INVX2_19/Y gnd NOR2X1_17/B vdd NAND3X1
XNAND3X1_92 INVX2_60/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_94/B vdd NAND3X1
XNOR2X1_70 NOR2X1_70/A NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_92 INVX2_81/A NOR2X1_93/B gnd NOR2X1_92/Y vdd NOR2X1
XNOR2X1_81 INVX2_89/A NOR2X1_82/B gnd NOR2X1_81/Y vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd ss_pad_o[5] vdd BUFX2
XNAND2X1_116 NAND3X1_258/Y NAND3X1_260/Y gnd INVX1_131/A vdd NAND2X1
XNAND2X1_127 OAI21X1_248/Y OAI21X1_250/Y gnd NOR2X1_72/B vdd NAND2X1
XNAND2X1_105 MUX2X1_10/Y BUFX4_63/Y gnd AOI21X1_42/B vdd NAND2X1
XNAND2X1_138 OAI21X1_273/Y OAI21X1_278/Y gnd OAI21X1_279/B vdd NAND2X1
XNAND2X1_3 BUFX4_90/Y wb_dat_i[26] gnd OAI21X1_5/C vdd NAND2X1
XNAND2X1_149 BUFX4_90/Y wb_dat_i[30] gnd OAI21X1_508/C vdd NAND2X1
XNOR2X1_160 INVX2_159/Y INVX2_154/A gnd NOR2X1_160/Y vdd NOR2X1
XOAI21X1_633 INVX4_10/A INVX8_20/Y MUX2X1_34/Y gnd OAI21X1_634/C vdd OAI21X1
XNOR2X1_193 INVX8_18/A NOR2X1_193/B gnd INVX1_152/A vdd NOR2X1
XOAI21X1_644 INVX1_121/Y BUFX4_19/Y OAI21X1_644/C gnd OAI21X1_644/Y vdd OAI21X1
XOAI21X1_600 INVX8_9/A INVX8_20/Y MUX2X1_28/Y gnd OAI21X1_601/C vdd OAI21X1
XOAI21X1_655 BUFX4_166/Y MUX2X1_39/Y OAI21X1_655/C gnd DFFSR_119/D vdd OAI21X1
XOAI21X1_666 BUFX4_234/Y OAI21X1_666/B BUFX4_45/Y gnd OAI22X1_118/D vdd OAI21X1
XOAI21X1_622 INVX1_156/Y INVX1_103/A BUFX4_165/Y gnd OAI21X1_623/B vdd OAI21X1
XOAI21X1_611 AND2X2_23/B INVX1_119/A BUFX4_161/Y gnd OAI21X1_612/B vdd OAI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNOR2X1_171 OR2X2_13/B NOR2X1_201/B gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_182 NOR2X1_202/B INVX8_19/Y gnd NOR2X1_182/Y vdd NOR2X1
XAOI21X1_8 INVX1_99/A BUFX4_114/Y AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XOAI21X1_699 INVX1_98/A NOR2X1_252/Y OAI21X1_699/C gnd OAI21X1_700/A vdd OAI21X1
XOAI21X1_688 BUFX4_157/Y OAI21X1_688/B OAI21X1_688/C gnd AOI22X1_87/C vdd OAI21X1
XOAI21X1_677 BUFX4_155/Y OR2X2_13/Y OAI21X1_677/C gnd AOI22X1_85/C vdd OAI21X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_73 INVX2_33/A gnd INVX1_73/Y vdd INVX1
XINVX1_51 INVX2_58/A gnd INVX1_51/Y vdd INVX1
XBUFX2_15 BUFX2_15/A gnd ss_pad_o[12] vdd BUFX2
XINVX1_62 INVX2_71/A gnd INVX1_62/Y vdd INVX1
XBUFX2_26 BUFX2_26/A gnd ss_pad_o[23] vdd BUFX2
XINVX1_40 INVX2_77/A gnd INVX1_40/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XBUFX2_37 DFFSR_66/Q gnd wb_dat_o[1] vdd BUFX2
XBUFX2_48 DFFSR_77/Q gnd wb_dat_o[12] vdd BUFX2
XBUFX2_59 DFFSR_88/Q gnd wb_dat_o[23] vdd BUFX2
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 MUX2X1_31/B BUFX4_114/Y OAI22X1_44/Y gnd NAND2X1_49/B vdd AOI21X1
XAOI21X1_27 AOI21X1_27/A AOI21X1_27/B NOR2X1_47/Y gnd DFFSR_114/D vdd AOI21X1
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B BUFX4_65/Y gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_49 AOI21X1_49/A AOI21X1_49/B INVX8_13/Y gnd AOI21X1_49/Y vdd AOI21X1
XFILL_26_4_0 gnd vdd FILL
XOAI22X1_57 OAI22X1_57/A NOR2X1_90/Y NOR2X1_91/Y OAI22X1_57/D gnd OAI22X1_57/Y vdd
+ OAI22X1
XOAI22X1_35 BUFX4_193/Y INVX2_5/Y INVX2_34/Y BUFX4_220/Y gnd NOR2X1_13/A vdd OAI22X1
XOAI22X1_46 OAI22X1_8/A INVX2_9/Y BUFX4_133/Y INVX1_63/Y gnd OAI22X1_46/Y vdd OAI22X1
XFILL_1_4_0 gnd vdd FILL
XOAI22X1_13 OAI22X1_7/A INVX1_31/Y INVX1_30/Y OAI22X1_7/D gnd NOR2X1_6/B vdd OAI22X1
XOAI22X1_24 INVX8_5/A INVX1_41/Y INVX8_2/A INVX2_30/Y gnd AOI21X1_8/C vdd OAI22X1
XOAI21X1_430 NOR2X1_169/Y MUX2X1_7/B BUFX4_230/Y gnd OAI21X1_430/Y vdd OAI21X1
XOAI21X1_474 NOR2X1_176/Y MUX2X1_5/A BUFX4_231/Y gnd OAI21X1_474/Y vdd OAI21X1
XOAI21X1_485 BUFX4_233/Y OAI21X1_485/B BUFX4_42/Y gnd OAI22X1_96/D vdd OAI21X1
XOAI21X1_441 BUFX4_55/Y BUFX4_125/Y NOR2X1_154/Y gnd NOR2X1_201/B vdd OAI21X1
XOAI21X1_463 INVX2_147/Y BUFX4_185/Y OAI21X1_624/C gnd OAI21X1_464/B vdd OAI21X1
XOAI21X1_452 BUFX4_229/Y OAI21X1_452/B INVX8_16/A gnd OAI22X1_90/D vdd OAI21X1
XOAI22X1_79 OAI22X1_79/A OAI22X1_79/B OAI22X1_79/C OAI22X1_79/D gnd OAI22X1_79/Y vdd
+ OAI22X1
XOAI21X1_496 INVX2_63/Y BUFX4_106/Y OAI21X1_573/C gnd OAI21X1_497/B vdd OAI21X1
XOAI22X1_68 OAI22X1_68/A OAI22X1_68/B OAI22X1_68/C OAI22X1_68/D gnd OAI22X1_68/Y vdd
+ OAI22X1
XFILL_9_5_0 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XOAI21X1_90 AND2X2_2/Y INVX2_29/Y OAI21X1_90/C gnd DFFSR_39/D vdd OAI21X1
XOAI21X1_260 AOI21X1_72/Y INVX2_151/Y INVX1_129/A gnd OAI21X1_260/Y vdd OAI21X1
XOAI21X1_271 NOR2X1_87/B MUX2X1_37/B BUFX4_37/Y gnd OAI22X1_56/A vdd OAI21X1
XOAI21X1_282 INVX1_20/A BUFX4_222/Y BUFX4_169/Y gnd OAI22X1_59/A vdd OAI21X1
XOAI21X1_293 INVX2_136/A NOR2X1_98/B BUFX4_80/Y gnd OAI22X1_63/D vdd OAI21X1
XFILL_29_3 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_23_2_0 gnd vdd FILL
XDFFSR_60 INVX2_36/A CLKBUF1_3/A DFFSR_2/R vdd DFFSR_60/D gnd vdd DFFSR
XDFFSR_82 DFFSR_82/Q DFFSR_82/CLK DFFSR_95/R vdd DFFSR_82/D gnd vdd DFFSR
XDFFSR_71 DFFSR_71/Q DFFSR_71/CLK DFFSR_3/R vdd DFFSR_71/D gnd vdd DFFSR
XDFFSR_93 DFFSR_93/Q DFFSR_93/CLK DFFSR_93/R vdd DFFSR_93/D gnd vdd DFFSR
XFILL_6_3_0 gnd vdd FILL
XFILL_15_7_1 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_132 NOR2X1_94/B gnd NOR2X1_74/B vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_110 MUX2X1_29/B gnd MUX2X1_30/B vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XAOI21X1_114 MUX2X1_4/A OAI21X1_386/B BUFX4_263/Y gnd OAI21X1_386/C vdd AOI21X1
XAOI21X1_103 AOI21X1_103/A NAND2X1_172/Y AND2X2_14/Y gnd OAI21X1_374/A vdd AOI21X1
XAOI21X1_125 BUFX4_263/Y OAI21X1_398/Y BUFX4_243/Y gnd AOI22X1_55/D vdd AOI21X1
XAOI21X1_158 NOR2X1_181/Y BUFX4_154/Y OAI21X1_489/Y gnd OAI22X1_98/C vdd AOI21X1
XAOI21X1_169 BUFX4_257/Y OAI21X1_520/Y BUFX4_5/Y gnd AOI22X1_70/D vdd AOI21X1
XAOI21X1_147 INVX2_123/Y OR2X2_12/Y BUFX4_255/Y gnd OAI21X1_454/C vdd AOI21X1
XAOI21X1_136 INVX2_105/Y OAI21X1_410/B BUFX4_254/Y gnd OAI21X1_410/C vdd AOI21X1
XNAND3X1_118 INVX2_75/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_119/C vdd NAND3X1
XNAND3X1_129 INVX2_91/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_130/C vdd NAND3X1
XNAND3X1_107 INVX2_68/Y BUFX4_76/Y BUFX4_57/Y gnd AOI21X1_36/A vdd NAND3X1
XFILL_30_5_1 gnd vdd FILL
XDFFSR_105 XNOR2X1_1/B CLKBUF1_5/A vdd DFFSR_115/S DFFSR_105/D gnd vdd DFFSR
XDFFSR_127 INVX1_92/A DFFSR_37/CLK BUFX4_14/Y vdd DFFSR_127/D gnd vdd DFFSR
XDFFSR_116 MUX2X1_43/B DFFSR_41/CLK BUFX4_18/Y vdd DFFSR_116/D gnd vdd DFFSR
XDFFSR_149 INVX2_95/A CLKBUF1_9/A BUFX4_18/Y vdd DFFSR_149/D gnd vdd DFFSR
XDFFSR_138 MUX2X1_29/B DFFSR_3/CLK BUFX4_13/Y vdd DFFSR_138/D gnd vdd DFFSR
XBUFX4_271 DFFSR_44/Q gnd OR2X2_6/B vdd BUFX4
XBUFX4_260 BUFX4_260/A gnd BUFX4_260/Y vdd BUFX4
XFILL_21_5_1 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_4_6_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd XOR2X1_5/B vdd NOR2X1
XNOR2X1_82 INVX2_90/A NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XFILL_19_1_0 gnd vdd FILL
XNAND3X1_60 BUFX4_200/Y NAND3X1_60/B BUFX4_130/Y gnd NAND3X1_60/Y vdd NAND3X1
XNAND3X1_71 wb_adr_i[2] wb_adr_i[3] INVX4_1/Y gnd INVX8_5/A vdd NAND3X1
XNAND3X1_93 INVX2_61/Y BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_94/C vdd NAND3X1
XNAND3X1_82 NAND3X1_82/A NAND3X1_82/B NAND3X1_82/C gnd DFFSR_91/D vdd NAND3X1
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XNOR2X1_93 INVX2_82/A NOR2X1_93/B gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd ss_pad_o[6] vdd BUFX2
XNAND2X1_117 AOI21X1_72/A AOI21X1_72/B gnd AOI21X1_66/A vdd NAND2X1
XNAND2X1_139 MUX2X1_1/A INVX4_8/A gnd OAI21X1_280/C vdd NAND2X1
XNAND2X1_128 BUFX4_181/Y OAI21X1_251/Y gnd OAI21X1_252/C vdd NAND2X1
XNAND2X1_106 MUX2X1_11/Y NOR2X1_66/B gnd AOI21X1_43/A vdd NAND2X1
XNAND2X1_4 BUFX4_92/Y wb_dat_i[27] gnd OAI21X1_7/C vdd NAND2X1
XNOR2X1_194 INVX4_11/Y INVX1_152/Y gnd NOR2X1_194/Y vdd NOR2X1
XNOR2X1_150 INVX2_157/Y INVX2_155/A gnd INVX1_142/A vdd NOR2X1
XNOR2X1_183 OR2X2_12/B INVX8_19/Y gnd NOR2X1_183/Y vdd NOR2X1
XNOR2X1_161 NOR2X1_71/A INVX1_138/Y gnd INVX1_139/A vdd NOR2X1
XNOR2X1_172 NOR2X1_202/B OR2X2_13/B gnd NOR2X1_172/Y vdd NOR2X1
XOAI21X1_634 MUX2X1_26/S MUX2X1_33/Y OAI21X1_634/C gnd DFFSR_128/D vdd OAI21X1
XOAI21X1_645 AND2X2_29/B INVX1_121/A BUFX4_166/Y gnd OAI21X1_646/B vdd OAI21X1
XAOI21X1_9 INVX1_121/A BUFX4_115/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_667 BUFX4_153/Y OAI21X1_667/B OAI21X1_667/C gnd AOI22X1_82/C vdd OAI21X1
XOAI21X1_678 INVX2_75/Y BUFX4_188/Y OAI21X1_697/C gnd OAI21X1_679/B vdd OAI21X1
XOAI21X1_623 NOR2X1_227/Y OAI21X1_623/B OAI21X1_623/C gnd DFFSR_133/D vdd OAI21X1
XOAI21X1_612 AND2X2_23/Y OAI21X1_612/B OAI21X1_612/C gnd DFFSR_136/D vdd OAI21X1
XOAI21X1_689 INVX2_74/Y BUFX4_189/Y OAI21X1_697/C gnd OAI21X1_689/Y vdd OAI21X1
XOAI21X1_656 BUFX4_127/Y INVX8_20/Y MUX2X1_42/Y gnd OAI21X1_657/C vdd OAI21X1
XOAI21X1_601 BUFX4_163/Y MUX2X1_27/Y OAI21X1_601/C gnd DFFSR_140/D vdd OAI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_52 INVX2_53/A gnd INVX1_52/Y vdd INVX1
XBUFX2_49 DFFSR_78/Q gnd wb_dat_o[13] vdd BUFX2
XBUFX2_16 BUFX2_16/A gnd ss_pad_o[13] vdd BUFX2
XINVX1_63 INVX2_70/A gnd INVX1_63/Y vdd INVX1
XBUFX2_38 DFFSR_67/Q gnd wb_dat_o[2] vdd BUFX2
XBUFX2_27 BUFX2_27/A gnd ss_pad_o[24] vdd BUFX2
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_41 INVX2_76/A gnd INVX1_41/Y vdd INVX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XAOI21X1_28 NOR2X1_62/A XOR2X1_5/B NOR2X1_60/A gnd NAND2X1_92/A vdd AOI21X1
XAOI21X1_17 INVX2_72/A BUFX4_68/Y OAI22X1_45/Y gnd NAND2X1_50/A vdd AOI21X1
XAOI21X1_39 AOI21X1_39/A AOI21X1_39/B BUFX4_81/Y gnd AOI21X1_39/Y vdd AOI21X1
XFILL_26_4_1 gnd vdd FILL
XOAI22X1_47 DFFSR_64/Q INVX1_64/Y OAI22X1_47/C INVX2_22/Y gnd DFFSR_63/D vdd OAI22X1
XOAI22X1_58 OAI22X1_58/A NOR2X1_92/Y NOR2X1_93/Y OAI22X1_58/D gnd OAI22X1_58/Y vdd
+ OAI22X1
XOAI22X1_36 INVX8_5/A INVX1_53/Y INVX8_2/A INVX2_21/Y gnd OAI22X1_36/Y vdd OAI22X1
XOAI22X1_25 OAI22X1_4/A INVX1_43/Y INVX1_42/Y INVX8_7/A gnd NOR2X1_10/B vdd OAI22X1
XOAI22X1_69 OAI22X1_69/A OAI22X1_69/B OAI22X1_69/C OAI22X1_69/D gnd OAI22X1_69/Y vdd
+ OAI22X1
XFILL_1_4_1 gnd vdd FILL
XOAI22X1_14 OAI22X1_8/A INVX2_14/Y INVX2_43/Y OAI22X1_8/D gnd NOR2X1_6/A vdd OAI22X1
XOAI21X1_431 MUX2X1_7/B BUFX4_88/Y OAI21X1_522/C gnd OAI21X1_432/B vdd OAI21X1
XOAI21X1_420 BUFX4_230/Y OAI21X1_420/B BUFX4_43/Y gnd OAI22X1_84/D vdd OAI21X1
XOAI21X1_475 MUX2X1_5/A BUFX4_26/Y OAI21X1_635/C gnd OAI21X1_476/B vdd OAI21X1
XOAI21X1_464 BUFX4_146/Y OAI21X1_464/B BUFX4_249/Y gnd AOI22X1_66/D vdd OAI21X1
XOAI21X1_453 BUFX4_54/Y BUFX4_126/Y NOR2X1_157/Y gnd OR2X2_12/B vdd OAI21X1
XOAI21X1_442 NOR2X1_171/Y INVX2_99/Y BUFX4_229/Y gnd OAI21X1_442/Y vdd OAI21X1
XOAI21X1_497 BUFX4_229/Y OAI21X1_497/B INVX8_16/A gnd OAI22X1_99/D vdd OAI21X1
XOAI21X1_486 NOR2X1_180/Y INVX2_114/Y BUFX4_234/Y gnd OAI21X1_486/Y vdd OAI21X1
XFILL_8_0_0 gnd vdd FILL
XFILL_9_5_1 gnd vdd FILL
XFILL_17_4_1 gnd vdd FILL
XOAI21X1_80 AND2X2_2/Y INVX2_24/Y OAI21X1_80/C gnd DFFSR_34/D vdd OAI21X1
XOAI21X1_91 INVX2_30/Y MUX2X1_47/S OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XOAI21X1_250 INVX1_131/Y AOI21X1_75/B AOI21X1_75/Y gnd OAI21X1_250/Y vdd OAI21X1
XOAI21X1_261 NOR2X1_87/B INVX1_104/A BUFX4_37/Y gnd OAI22X1_52/A vdd OAI21X1
XOAI21X1_283 INVX2_145/A NOR2X1_98/B BUFX4_79/Y gnd OAI22X1_59/D vdd OAI21X1
XOAI21X1_294 NOR2X1_96/B INVX1_118/A BUFX4_39/Y gnd OAI22X1_64/A vdd OAI21X1
XOAI21X1_272 NOR2X1_78/B INVX1_105/A BUFX4_32/Y gnd OAI22X1_56/D vdd OAI21X1
XFILL_23_2_1 gnd vdd FILL
XDFFSR_50 INVX2_42/A CLKBUF1_3/Y DFFSR_63/R vdd DFFSR_50/D gnd vdd DFFSR
XDFFSR_94 DFFSR_94/Q DFFSR_4/CLK DFFSR_2/R vdd DFFSR_94/D gnd vdd DFFSR
XDFFSR_83 DFFSR_83/Q DFFSR_83/CLK DFFSR_95/R vdd DFFSR_83/D gnd vdd DFFSR
XDFFSR_72 DFFSR_72/Q DFFSR_87/CLK DFFSR_9/R vdd DFFSR_72/D gnd vdd DFFSR
XDFFSR_61 INVX2_37/A DFFSR_91/CLK DFFSR_9/R vdd DFFSR_61/D gnd vdd DFFSR
XFILL_6_3_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_133 XOR2X1_6/Y gnd NOR2X1_94/A vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_144 BUFX4_35/Y gnd INVX1_144/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_111 MUX2X1_35/B gnd MUX2X1_36/B vdd INVX1
XAOI21X1_115 BUFX4_263/Y OAI21X1_387/Y BUFX4_243/Y gnd AOI22X1_51/D vdd AOI21X1
XAOI21X1_137 NOR2X1_165/Y BUFX4_154/Y OAI21X1_414/Y gnd OAI22X1_83/C vdd AOI21X1
XAOI21X1_104 INVX2_92/Y OAI21X1_375/B BUFX4_266/Y gnd OAI21X1_375/C vdd AOI21X1
XAOI21X1_148 INVX2_91/Y OAI21X1_458/B BUFX4_255/Y gnd OAI21X1_458/C vdd AOI21X1
XAOI21X1_126 INVX2_133/Y OAI21X1_399/B BUFX4_262/Y gnd OAI21X1_399/C vdd AOI21X1
XAOI21X1_159 INVX2_135/Y OAI21X1_492/B BUFX4_254/Y gnd OAI21X1_492/C vdd AOI21X1
XNAND3X1_108 INVX2_69/Y BUFX4_48/Y BUFX4_138/Y gnd AOI21X1_36/B vdd NAND3X1
XNAND3X1_119 BUFX4_62/Y NAND3X1_119/B NAND3X1_119/C gnd AOI21X1_39/B vdd NAND3X1
XDFFSR_106 NOR2X1_27/B DFFSR_1/CLK vdd DFFSR_99/R DFFSR_106/D gnd vdd DFFSR
XDFFSR_128 MUX2X1_33/B DFFSR_98/CLK BUFX4_14/Y vdd DFFSR_128/D gnd vdd DFFSR
XDFFSR_117 INVX1_104/A CLKBUF1_25/Y BUFX4_18/Y vdd DFFSR_117/D gnd vdd DFFSR
XDFFSR_139 INVX1_98/A CLKBUF1_7/Y BUFX4_12/Y vdd DFFSR_139/D gnd vdd DFFSR
XBUFX4_272 DFFSR_44/Q gnd BUFX4_272/Y vdd BUFX4
XBUFX4_250 BUFX4_250/A gnd BUFX4_250/Y vdd BUFX4
XBUFX4_261 BUFX4_268/A gnd BUFX4_261/Y vdd BUFX4
XFILL_20_0_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 OAI21X1_91/Y AND2X2_3/B INVX8_2/Y gnd OAI21X1_92/C vdd NAND3X1
XNOR2X1_50 XOR2X1_3/A OR2X2_4/Y gnd INVX1_81/A vdd NOR2X1
XNOR2X1_61 INVX2_52/A INVX2_48/Y gnd NOR2X1_62/B vdd NOR2X1
XNAND3X1_83 NAND3X1_83/A NAND3X1_83/B NAND3X1_83/C gnd DFFSR_92/D vdd NAND3X1
XNOR2X1_72 NOR2X1_85/A NOR2X1_72/B gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_83 INVX2_87/A NOR2X1_84/B gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_94 NOR2X1_94/A NOR2X1_94/B gnd NOR2X1_94/Y vdd NOR2X1
XNAND3X1_61 BUFX4_202/Y NAND3X1_61/B AND2X2_3/A gnd NAND3X1_61/Y vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNAND3X1_72 NAND3X1_72/A AOI22X1_2/Y AOI22X1_1/Y gnd DFFSR_81/D vdd NAND3X1
XNAND3X1_94 BUFX4_206/Y NAND3X1_94/B NAND3X1_94/C gnd NAND3X1_94/Y vdd NAND3X1
XNAND2X1_107 MUX2X1_12/Y BUFX4_63/Y gnd AOI21X1_43/B vdd NAND2X1
XNAND2X1_118 INVX2_48/Y NOR3X1_5/Y gnd NAND3X1_263/B vdd NAND2X1
XNAND2X1_129 BUFX4_183/Y OAI21X1_254/Y gnd NAND2X1_132/A vdd NAND2X1
XNAND2X1_5 BUFX4_87/Y wb_dat_i[28] gnd OAI21X1_9/C vdd NAND2X1
XNOR2X1_151 INVX2_158/Y INVX2_155/A gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_195 BUFX4_253/Y NOR2X1_195/B gnd NOR2X1_195/Y vdd NOR2X1
XNOR2X1_184 INVX1_147/A INVX8_19/Y gnd NOR2X1_184/Y vdd NOR2X1
XNOR2X1_173 NOR2X1_71/A INVX1_149/Y gnd INVX8_19/A vdd NOR2X1
XNOR2X1_162 INVX1_140/Y INVX1_139/Y gnd INVX1_141/A vdd NOR2X1
XNOR2X1_140 INVX2_116/A BUFX4_179/Y gnd OAI22X1_81/C vdd NOR2X1
XOAI21X1_635 MUX2X1_3/A BUFX4_24/Y OAI21X1_635/C gnd OAI21X1_635/Y vdd OAI21X1
XOAI21X1_646 AND2X2_29/Y OAI21X1_646/B OAI21X1_646/C gnd DFFSR_124/D vdd OAI21X1
XOAI21X1_668 INVX2_72/Y BUFX4_21/Y OAI21X1_694/C gnd OAI21X1_668/Y vdd OAI21X1
XOAI21X1_679 BUFX4_145/Y OAI21X1_679/B BUFX4_244/Y gnd AOI22X1_85/D vdd OAI21X1
XOAI21X1_624 INVX1_122/Y BUFX4_185/Y OAI21X1_624/C gnd OAI21X1_624/Y vdd OAI21X1
XOAI21X1_657 BUFX4_161/Y MUX2X1_41/Y OAI21X1_657/C gnd DFFSR_118/D vdd OAI21X1
XOAI21X1_602 BUFX4_127/Y INVX8_22/Y AND2X2_18/A gnd NOR2X1_237/B vdd OAI21X1
XOAI21X1_613 INVX1_94/Y BUFX4_189/Y OAI21X1_613/C gnd OAI21X1_613/Y vdd OAI21X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XBUFX2_39 DFFSR_68/Q gnd wb_dat_o[3] vdd BUFX2
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_75 INVX1_75/A gnd NOR3X1_2/B vdd INVX1
XINVX1_53 INVX2_56/A gnd INVX1_53/Y vdd INVX1
XBUFX2_28 BUFX2_28/A gnd ss_pad_o[25] vdd BUFX2
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XBUFX2_17 BUFX2_17/A gnd ss_pad_o[14] vdd BUFX2
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_29 NAND2X1_92/A NAND3X1_91/Y INVX1_90/Y gnd AOI21X1_29/Y vdd AOI21X1
XAOI21X1_18 INVX1_97/A BUFX4_114/Y OAI22X1_46/Y gnd NAND2X1_50/B vdd AOI21X1
XOAI22X1_48 OR2X2_3/A OAI22X1_49/A OAI22X1_49/C OAI22X1_48/D gnd DFFSR_97/D vdd OAI22X1
XOAI21X1_432 BUFX4_230/Y OAI21X1_432/B BUFX4_44/Y gnd OAI22X1_87/D vdd OAI21X1
XOAI22X1_37 NOR2X1_18/B INVX1_55/Y INVX1_54/Y BUFX4_134/Y gnd NOR2X1_14/B vdd OAI22X1
XOAI21X1_421 BUFX4_52/Y BUFX4_125/Y NOR2X1_149/Y gnd NOR2X1_193/B vdd OAI21X1
XOAI22X1_26 OAI22X1_5/A INVX2_2/Y INVX2_31/Y INVX8_4/A gnd NOR2X1_10/A vdd OAI22X1
XOAI21X1_410 BUFX4_158/Y OAI21X1_410/B OAI21X1_410/C gnd AOI22X1_61/C vdd OAI21X1
XOAI22X1_59 OAI22X1_59/A NOR2X1_95/Y NOR2X1_96/Y OAI22X1_59/D gnd OAI22X1_59/Y vdd
+ OAI22X1
XOAI22X1_15 INVX8_5/A INVX1_32/Y INVX8_2/A INVX2_27/Y gnd AOI21X1_5/C vdd OAI22X1
XOAI21X1_476 BUFX4_231/Y OAI21X1_476/B BUFX4_43/Y gnd OAI22X1_93/D vdd OAI21X1
XOAI21X1_454 BUFX4_158/Y OR2X2_12/Y OAI21X1_454/C gnd AOI22X1_64/C vdd OAI21X1
XOAI21X1_498 NOR2X1_183/Y INVX2_126/Y BUFX4_229/Y gnd OAI21X1_498/Y vdd OAI21X1
XOAI21X1_443 INVX2_99/Y BUFX4_187/Y OAI21X1_605/C gnd OAI21X1_444/B vdd OAI21X1
XOAI21X1_465 BUFX4_155/Y OAI21X1_465/B OAI21X1_465/C gnd AOI22X1_67/C vdd OAI21X1
XOAI21X1_487 INVX2_114/Y BUFX4_111/Y OAI21X1_567/C gnd OAI21X1_488/B vdd OAI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_70 AND2X2_2/Y INVX2_21/Y OAI21X1_70/C gnd DFFSR_44/D vdd OAI21X1
XOAI21X1_81 INVX2_25/Y MUX2X1_43/S OAI21X1_81/C gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_92 AND2X2_2/Y INVX2_30/Y OAI21X1_92/C gnd DFFSR_40/D vdd OAI21X1
XFILL_27_7_0 gnd vdd FILL
XFILL_2_7_0 gnd vdd FILL
XOAI21X1_240 NOR3X1_6/C NOR3X1_6/B NOR3X1_6/A gnd OAI21X1_241/C vdd OAI21X1
XOAI21X1_251 NOR2X1_256/B INVX4_8/A OAI21X1_251/C gnd OAI21X1_251/Y vdd OAI21X1
XOAI21X1_273 OAI22X1_55/Y OAI22X1_56/Y NOR2X1_85/Y gnd OAI21X1_273/Y vdd OAI21X1
XOAI21X1_262 NOR2X1_78/B INVX1_103/A BUFX4_32/Y gnd OAI22X1_52/D vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_295 BUFX4_176/Y INVX1_119/A BUFX4_35/Y gnd OAI22X1_64/D vdd OAI21X1
XOAI21X1_284 NOR2X1_96/B MUX2X1_43/B BUFX4_39/Y gnd OAI22X1_60/A vdd OAI21X1
XFILL_18_7_0 gnd vdd FILL
XDFFSR_40 INVX2_30/A DFFSR_55/CLK DFFSR_63/R vdd DFFSR_40/D gnd vdd DFFSR
XDFFSR_62 INVX2_38/A DFFSR_2/CLK DFFSR_2/R vdd DFFSR_62/D gnd vdd DFFSR
XDFFSR_95 DFFSR_95/Q DFFSR_5/CLK DFFSR_95/R vdd DFFSR_95/D gnd vdd DFFSR
XDFFSR_73 DFFSR_73/Q DFFSR_88/CLK DFFSR_3/R vdd DFFSR_73/D gnd vdd DFFSR
XDFFSR_84 DFFSR_84/Q DFFSR_9/CLK DFFSR_3/R vdd DFFSR_84/D gnd vdd DFFSR
XDFFSR_51 INVX2_43/A DFFSR_96/CLK DFFSR_9/R vdd DFFSR_51/D gnd vdd DFFSR
XCLKBUF1_60 wb_clk_i gnd CLKBUF1_60/Y vdd CLKBUF1
XINVX1_134 NOR3X1_9/A gnd INVX1_134/Y vdd INVX1
XINVX1_101 INVX1_101/A gnd MUX2X1_12/A vdd INVX1
XINVX1_112 MUX2X1_23/B gnd MUX2X1_24/B vdd INVX1
XINVX1_123 MUX2X1_43/B gnd MUX2X1_44/B vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XAOI21X1_138 NOR2X1_166/Y BUFX4_152/Y OAI21X1_418/Y gnd OAI22X1_84/C vdd AOI21X1
XAOI21X1_105 BUFX4_266/Y OAI21X1_376/Y BUFX4_249/Y gnd AOI22X1_47/D vdd AOI21X1
XAOI21X1_149 INVX2_147/Y OAI21X1_462/B BUFX4_254/Y gnd OAI21X1_462/C vdd AOI21X1
XAOI21X1_127 BUFX4_261/Y OAI21X1_400/Y BUFX4_245/Y gnd AOI22X1_56/D vdd AOI21X1
XAOI21X1_116 INVX2_118/Y INVX1_143/Y BUFX4_268/Y gnd AOI21X1_117/A vdd AOI21X1
XFILL_24_5_0 gnd vdd FILL
XNAND3X1_109 INVX1_97/Y BUFX4_48/Y BUFX4_138/Y gnd AOI21X1_37/A vdd NAND3X1
XFILL_7_6_0 gnd vdd FILL
XDFFSR_107 NOR2X1_26/B DFFSR_2/CLK vdd DFFSR_108/S DFFSR_107/D gnd vdd DFFSR
XFILL_15_5_0 gnd vdd FILL
XDFFSR_129 INVX1_101/A CLKBUF1_37/Y BUFX4_18/Y vdd DFFSR_129/D gnd vdd DFFSR
XDFFSR_118 MUX2X1_41/B DFFSR_88/CLK BUFX4_13/Y vdd DFFSR_118/D gnd vdd DFFSR
XBUFX4_240 BUFX4_242/A gnd NOR2X1_18/B vdd BUFX4
XBUFX4_251 BUFX4_255/A gnd BUFX4_251/Y vdd BUFX4
XBUFX4_262 BUFX4_268/A gnd BUFX4_262/Y vdd BUFX4
XBUFX4_273 BUFX4_277/A gnd INVX8_14/A vdd BUFX4
XNAND3X1_84 NAND3X1_84/A NAND3X1_84/B NAND3X1_84/C gnd DFFSR_93/D vdd NAND3X1
XNAND3X1_40 OAI21X1_73/Y AND2X2_3/B INVX8_2/Y gnd OAI21X1_74/C vdd NAND3X1
XNAND3X1_51 wb_adr_i[4] wb_adr_i[2] INVX2_19/Y gnd BUFX4_220/A vdd NAND3X1
XNAND3X1_73 NAND3X1_73/A AOI22X1_4/Y AOI22X1_3/Y gnd DFFSR_82/D vdd NAND3X1
XNAND3X1_62 BUFX4_199/Y NAND3X1_62/B BUFX4_129/Y gnd NAND3X1_62/Y vdd NAND3X1
XNOR2X1_40 NOR3X1_1/A NOR3X1_1/C gnd NOR2X1_43/B vdd NOR2X1
XNOR2X1_51 NOR2X1_51/A INVX1_81/Y gnd OR2X2_3/B vdd NOR2X1
XNOR2X1_73 OR2X2_8/B NOR2X1_73/B gnd XOR2X1_6/B vdd NOR2X1
XNOR2X1_84 INVX2_88/A NOR2X1_84/B gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_62 NOR2X1_62/A NOR2X1_62/B gnd XOR2X1_4/B vdd NOR2X1
XNOR2X1_95 INVX1_19/A NOR2X1_96/B gnd NOR2X1_95/Y vdd NOR2X1
XNAND3X1_95 INVX1_94/Y BUFX4_50/Y BUFX4_136/Y gnd NAND3X1_97/B vdd NAND3X1
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_119 INVX2_48/A NOR3X1_5/Y gnd NAND3X1_264/B vdd NAND2X1
XNAND2X1_108 MUX2X1_13/Y NOR2X1_66/B gnd NAND3X1_212/B vdd NAND2X1
XNAND2X1_6 BUFX4_89/Y wb_dat_i[29] gnd NAND2X1_6/Y vdd NAND2X1
XNOR2X1_196 INVX8_18/A NOR2X1_196/B gnd INVX1_153/A vdd NOR2X1
XFILL_21_3_0 gnd vdd FILL
XNOR2X1_174 INVX8_19/Y NOR2X1_189/B gnd NOR2X1_174/Y vdd NOR2X1
XNOR2X1_152 INVX2_159/Y INVX2_155/A gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_130 INVX2_123/A NOR2X1_98/B gnd OAI22X1_76/B vdd NOR2X1
XOAI21X1_603 BUFX4_124/Y INVX8_20/Y MUX2X1_30/Y gnd OAI21X1_604/C vdd OAI21X1
XNOR2X1_185 BUFX4_127/Y INVX8_20/Y gnd BUFX4_7/A vdd NOR2X1
XNOR2X1_163 INVX1_142/Y INVX1_139/Y gnd INVX1_143/A vdd NOR2X1
XOAI21X1_614 BUFX4_121/Y INVX8_22/Y AND2X2_20/A gnd NOR2X1_240/B vdd OAI21X1
XNOR2X1_141 INVX1_49/A BUFX4_179/Y gnd OAI22X1_81/B vdd NOR2X1
XOAI21X1_636 AND2X2_26/B INVX1_92/A BUFX4_162/Y gnd OAI21X1_637/B vdd OAI21X1
XOAI21X1_658 INVX1_104/Y BUFX4_106/Y OAI21X1_658/C gnd OAI21X1_658/Y vdd OAI21X1
XOAI21X1_625 BUFX4_127/Y INVX8_22/Y NOR2X1_205/Y gnd NOR2X1_243/B vdd OAI21X1
XOAI21X1_669 BUFX4_155/Y OAI21X1_669/B OAI21X1_669/C gnd AOI22X1_83/C vdd OAI21X1
XOAI21X1_647 BUFX4_124/Y INVX8_20/Y MUX2X1_36/Y gnd OAI21X1_648/C vdd OAI21X1
XINVX1_65 XOR2X1_1/B gnd INVX1_65/Y vdd INVX1
XINVX1_76 NOR3X1_2/A gnd INVX1_76/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_21 INVX2_96/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XFILL_29_4_0 gnd vdd FILL
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XBUFX2_29 BUFX2_29/A gnd ss_pad_o[26] vdd BUFX2
XFILL_4_4_0 gnd vdd FILL
XBUFX2_18 BUFX2_18/A gnd ss_pad_o[15] vdd BUFX2
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND3X1_270 AOI21X1_72/A NOR3X1_7/C AOI21X1_72/B gnd NAND3X1_271/B vdd NAND3X1
XAOI21X1_19 INVX1_17/A OR2X2_1/A OR2X2_1/B gnd OAI22X1_48/D vdd AOI21X1
XOAI22X1_49 OAI22X1_49/A OAI22X1_49/B OAI22X1_49/C OR2X2_3/A gnd DFFSR_98/D vdd OAI22X1
XOAI21X1_422 NOR2X1_167/Y MUX2X1_5/B BUFX4_231/Y gnd OAI21X1_422/Y vdd OAI21X1
XOAI22X1_38 BUFX4_193/Y INVX2_6/Y INVX2_35/Y BUFX4_220/Y gnd NOR2X1_14/A vdd OAI22X1
XOAI22X1_16 BUFX4_193/Y INVX2_15/Y INVX2_44/Y BUFX4_220/Y gnd NOR2X1_7/A vdd OAI22X1
XOAI21X1_433 BUFX4_52/Y BUFX4_125/Y NOR2X1_152/Y gnd NOR2X1_198/B vdd OAI21X1
XOAI22X1_27 INVX8_5/A INVX1_44/Y INVX8_2/A INVX1_17/Y gnd AOI21X1_9/C vdd OAI22X1
XOAI21X1_455 INVX2_123/Y BUFX4_190/Y OAI21X1_617/C gnd OAI21X1_456/B vdd OAI21X1
XOAI21X1_411 INVX2_105/Y BUFX4_90/Y OAI21X1_508/C gnd OAI21X1_412/B vdd OAI21X1
XOAI21X1_444 BUFX4_229/Y OAI21X1_444/B INVX8_16/A gnd OAI22X1_89/D vdd OAI21X1
XOAI21X1_400 INVX2_133/Y MUX2X1_37/S OAI21X1_651/C gnd OAI21X1_400/Y vdd OAI21X1
XOAI21X1_466 INVX2_108/Y BUFX4_23/Y OAI21X1_548/C gnd OAI21X1_467/B vdd OAI21X1
XOAI21X1_477 NOR2X1_177/Y INVX2_120/Y BUFX4_232/Y gnd OAI21X1_477/Y vdd OAI21X1
XOAI21X1_499 INVX2_126/Y MUX2X1_43/S OAI21X1_575/C gnd OAI21X1_500/B vdd OAI21X1
XOAI21X1_488 BUFX4_234/Y OAI21X1_488/B BUFX4_45/Y gnd OAI22X1_97/D vdd OAI21X1
XOAI21X1_71 INVX2_22/Y BUFX4_22/Y OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_93 INVX2_31/Y BUFX4_25/Y OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_60 BUFX4_101/Y INVX2_15/Y OAI21X1_60/C gnd DFFSR_6/D vdd OAI21X1
XOAI21X1_82 AND2X2_2/Y INVX2_25/Y OAI21X1_82/C gnd DFFSR_35/D vdd OAI21X1
XFILL_27_7_1 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XFILL_2_7_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_241 NOR3X1_7/A INVX2_151/A OAI21X1_241/C gnd AOI21X1_66/C vdd OAI21X1
XOAI21X1_252 XNOR2X1_12/Y BUFX4_181/Y OAI21X1_252/C gnd NOR2X1_85/A vdd OAI21X1
XOAI21X1_274 INVX2_83/A NOR2X1_93/B BUFX4_168/Y gnd OAI22X1_57/A vdd OAI21X1
XOAI21X1_263 OAI22X1_51/Y OAI22X1_52/Y INVX2_154/Y gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_285 BUFX4_176/Y INVX1_122/A BUFX4_35/Y gnd OAI22X1_60/D vdd OAI21X1
XOAI21X1_296 OAI22X1_63/Y OAI22X1_64/Y NOR2X1_85/Y gnd OAI21X1_296/Y vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XOAI21X1_230 AOI21X1_57/Y AOI21X1_58/Y INVX4_5/A gnd AOI21X1_59/B vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XFILL_18_7_1 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XDFFSR_30 INVX1_6/A DFFSR_30/CLK DFFSR_3/R vdd DFFSR_30/D gnd vdd DFFSR
XDFFSR_74 DFFSR_74/Q CLKBUF1_3/A DFFSR_93/R vdd DFFSR_74/D gnd vdd DFFSR
XDFFSR_41 INVX1_17/A DFFSR_41/CLK DFFSR_93/R vdd DFFSR_41/D gnd vdd DFFSR
XDFFSR_63 INVX1_64/A DFFSR_93/CLK DFFSR_63/R vdd DFFSR_63/D gnd vdd DFFSR
XDFFSR_52 INVX2_44/A DFFSR_7/CLK DFFSR_63/R vdd DFFSR_52/D gnd vdd DFFSR
XDFFSR_85 DFFSR_85/Q DFFSR_85/CLK DFFSR_95/R vdd DFFSR_85/D gnd vdd DFFSR
XDFFSR_96 DFFSR_96/Q DFFSR_96/CLK DFFSR_96/R vdd DFFSR_96/D gnd vdd DFFSR
XCLKBUF1_61 wb_clk_i gnd CLKBUF1_61/Y vdd CLKBUF1
XCLKBUF1_50 CLKBUF1_57/Y gnd DFFSR_96/CLK vdd CLKBUF1
XINVX1_124 OR2X2_7/A gnd INVX1_124/Y vdd INVX1
XINVX1_135 NOR2X1_72/B gnd NOR2X1_85/B vdd INVX1
XINVX1_102 MUX2X1_19/B gnd MUX2X1_20/B vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XAOI21X1_139 NOR2X1_167/Y BUFX4_154/Y OAI21X1_422/Y gnd OAI22X1_85/C vdd AOI21X1
XAOI21X1_106 INVX2_145/Y OAI21X1_377/B BUFX4_266/Y gnd OAI21X1_377/C vdd AOI21X1
XAOI21X1_128 INVX2_64/Y OAI21X1_401/B BUFX4_261/Y gnd OAI21X1_401/C vdd AOI21X1
XAOI21X1_117 AOI21X1_117/A NAND2X1_186/Y AND2X2_16/Y gnd OAI21X1_390/A vdd AOI21X1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XINVX4_10 INVX4_10/A gnd INVX4_10/Y vdd INVX4
XFILL_6_1_0 gnd vdd FILL
XFILL_7_6_1 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XDFFSR_108 NOR3X1_1/B DFFSR_93/CLK vdd DFFSR_108/S DFFSR_108/D gnd vdd DFFSR
XFILL_14_0_0 gnd vdd FILL
XDFFSR_119 INVX1_95/A CLKBUF1_6/A BUFX4_11/Y vdd DFFSR_119/D gnd vdd DFFSR
XBUFX4_230 INVX8_18/Y gnd BUFX4_230/Y vdd BUFX4
XBUFX4_263 BUFX4_268/A gnd BUFX4_263/Y vdd BUFX4
XBUFX4_252 BUFX4_255/A gnd INVX8_18/A vdd BUFX4
XBUFX4_241 BUFX4_242/A gnd OAI22X1_4/A vdd BUFX4
XBUFX4_274 BUFX4_277/A gnd MUX2X1_48/A vdd BUFX4
XNOR2X1_30 INVX2_33/A INVX2_34/A gnd NOR2X1_30/Y vdd NOR2X1
XNAND3X1_41 OAI21X1_75/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_76/C vdd NAND3X1
XNAND3X1_52 BUFX4_202/Y OAI21X1_93/Y BUFX4_131/Y gnd OAI21X1_94/C vdd NAND3X1
XNAND3X1_63 BUFX4_200/Y NAND3X1_63/B BUFX4_130/Y gnd NAND3X1_63/Y vdd NAND3X1
XNAND3X1_85 NAND3X1_85/A NAND3X1_85/B NAND3X1_85/C gnd DFFSR_94/D vdd NAND3X1
XNAND3X1_30 AND2X2_3/B OAI21X1_55/Y BUFX4_97/Y gnd OAI21X1_56/C vdd NAND3X1
XNAND3X1_74 NAND3X1_74/A AOI22X1_6/Y AOI22X1_5/Y gnd DFFSR_83/D vdd NAND3X1
XNAND3X1_96 INVX2_62/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_97/C vdd NAND3X1
XNOR2X1_41 INVX1_70/A NOR3X1_1/C gnd XNOR2X1_1/A vdd NOR2X1
XNOR2X1_52 MUX2X1_1/Y OR2X2_3/B gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_63 XOR2X1_3/Y NOR2X1_64/B gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A NOR2X1_85/B gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_94/A NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_109 MUX2X1_14/Y BUFX4_66/Y gnd NAND3X1_212/C vdd NAND2X1
XNAND2X1_7 BUFX4_91/Y wb_dat_i[30] gnd NAND2X1_7/Y vdd NAND2X1
XNOR2X1_142 INVX2_117/A NOR2X1_79/B gnd OAI22X1_82/B vdd NOR2X1
XNOR2X1_131 INVX1_24/A BUFX4_222/Y gnd OAI22X1_76/C vdd NOR2X1
XNOR2X1_120 INVX2_74/A BUFX4_176/Y gnd OAI22X1_71/C vdd NOR2X1
XNOR2X1_197 INVX4_11/Y INVX1_153/Y gnd NOR2X1_197/Y vdd NOR2X1
XNOR2X1_175 INVX8_19/Y NOR2X1_191/B gnd NOR2X1_175/Y vdd NOR2X1
XOAI21X1_637 AND2X2_26/Y OAI21X1_637/B OAI21X1_637/C gnd DFFSR_127/D vdd OAI21X1
XFILL_21_3_1 gnd vdd FILL
XNOR2X1_153 INVX2_157/Y INVX2_160/Y gnd NOR2X1_153/Y vdd NOR2X1
XOAI21X1_626 INVX1_122/A NOR2X1_228/Y OAI21X1_626/C gnd OAI21X1_627/A vdd OAI21X1
XOAI21X1_604 BUFX4_161/Y MUX2X1_29/Y OAI21X1_604/C gnd DFFSR_138/D vdd OAI21X1
XNOR2X1_164 NOR2X1_98/B INVX1_144/Y gnd INVX8_17/A vdd NOR2X1
XOAI21X1_648 BUFX4_163/Y MUX2X1_35/Y OAI21X1_648/C gnd DFFSR_122/D vdd OAI21X1
XOAI21X1_615 INVX1_94/A NOR2X1_224/Y OAI21X1_615/C gnd OAI21X1_616/A vdd OAI21X1
XNOR2X1_186 BUFX4_179/Y NOR2X1_71/B gnd INVX4_11/A vdd NOR2X1
XOAI21X1_659 INVX1_157/Y INVX1_104/A BUFX4_166/Y gnd OAI21X1_660/B vdd OAI21X1
XFILL_29_4_1 gnd vdd FILL
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_77 NOR3X1_3/A gnd INVX1_77/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_66 INVX2_38/A gnd INVX1_66/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_22 INVX2_95/A gnd INVX1_22/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd ss_pad_o[16] vdd BUFX2
XFILL_12_3_1 gnd vdd FILL
XNAND3X1_260 INVX4_6/Y OAI21X1_237/Y NAND3X1_260/C gnd NAND3X1_260/Y vdd NAND3X1
XNAND3X1_271 BUFX4_272/Y NAND3X1_271/B NAND3X1_272/C gnd AND2X2_13/A vdd NAND3X1
XOAI22X1_28 NOR2X1_18/B INVX1_46/Y INVX1_45/Y BUFX4_134/Y gnd NOR2X1_11/B vdd OAI22X1
XOAI22X1_39 INVX8_5/A INVX1_56/Y INVX8_2/A INVX2_22/Y gnd OAI22X1_39/Y vdd OAI22X1
XOAI22X1_17 OAI22X1_4/A INVX1_34/Y INVX1_33/Y INVX8_7/A gnd NOR2X1_7/B vdd OAI22X1
XOAI21X1_423 MUX2X1_5/B BUFX4_86/Y OAI21X1_590/C gnd OAI21X1_424/B vdd OAI21X1
XOAI21X1_456 BUFX4_143/Y OAI21X1_456/B BUFX4_249/Y gnd AOI22X1_64/D vdd OAI21X1
XOAI21X1_489 NOR2X1_181/Y INVX2_102/Y BUFX4_232/Y gnd OAI21X1_489/Y vdd OAI21X1
XOAI21X1_434 NOR2X1_170/Y INVX2_141/Y BUFX4_232/Y gnd OAI21X1_434/Y vdd OAI21X1
XOAI21X1_478 INVX2_120/Y BUFX4_19/Y OAI21X1_638/C gnd OAI21X1_479/B vdd OAI21X1
XOAI21X1_412 BUFX4_145/Y OAI21X1_412/B BUFX4_244/Y gnd AOI22X1_61/D vdd OAI21X1
XOAI21X1_445 BUFX4_54/Y BUFX4_126/Y NOR2X1_155/Y gnd INVX1_146/A vdd OAI21X1
XOAI21X1_401 BUFX4_155/Y OAI21X1_401/B OAI21X1_401/C gnd AOI22X1_57/C vdd OAI21X1
XOAI21X1_467 BUFX4_144/Y OAI21X1_467/B BUFX4_245/Y gnd AOI22X1_67/D vdd OAI21X1
XOAI21X1_72 AND2X2_2/Y INVX2_22/Y OAI21X1_72/C gnd DFFSR_45/D vdd OAI21X1
XOAI21X1_94 AND2X2_3/Y INVX2_31/Y OAI21X1_94/C gnd DFFSR_55/D vdd OAI21X1
XOAI21X1_83 INVX2_26/Y BUFX4_108/Y OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_61 INVX2_16/Y MUX2X1_37/S OAI21X1_89/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_50 OAI21X1_8/A INVX2_10/Y OAI21X1_50/C gnd DFFSR_1/D vdd OAI21X1
XFILL_26_2_1 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_242 AND2X2_8/Y NOR2X1_54/A INVX4_8/A gnd AOI21X1_67/B vdd OAI21X1
XOAI21X1_253 AND2X2_8/Y NOR2X1_54/A INVX4_8/Y gnd OAI21X1_254/C vdd OAI21X1
XOAI21X1_220 MUX2X1_25/B MUX2X1_6/S OAI21X1_220/C gnd AND2X2_11/B vdd OAI21X1
XOAI21X1_275 INVX2_84/A NOR2X1_93/B BUFX4_77/Y gnd OAI22X1_57/D vdd OAI21X1
XOAI21X1_264 INVX2_85/A NOR2X1_84/B BUFX4_168/Y gnd OAI22X1_53/A vdd OAI21X1
XOAI21X1_231 AOI21X1_59/Y AOI21X1_54/Y INVX1_86/A gnd OAI21X1_231/Y vdd OAI21X1
XOAI21X1_297 INVX1_44/A NOR2X1_88/B BUFX4_168/Y gnd OAI22X1_65/A vdd OAI21X1
XAND2X2_20 AND2X2_20/A INVX4_11/A gnd AND2X2_20/Y vdd AND2X2
XOAI21X1_286 OAI22X1_59/Y OAI22X1_60/Y INVX2_154/Y gnd OAI21X1_286/Y vdd OAI21X1
XFILL_9_3_1 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XDFFSR_42 INVX4_8/A DFFSR_57/CLK DFFSR_93/R vdd DFFSR_42/D gnd vdd DFFSR
XDFFSR_53 INVX2_45/A DFFSR_8/CLK DFFSR_63/R vdd DFFSR_53/D gnd vdd DFFSR
XDFFSR_64 DFFSR_64/Q CLKBUF1_5/Y DFFSR_2/R vdd DFFSR_64/D gnd vdd DFFSR
XDFFSR_31 INVX1_7/A DFFSR_91/CLK DFFSR_96/R vdd DFFSR_31/D gnd vdd DFFSR
XDFFSR_20 INVX1_12/A DFFSR_5/CLK DFFSR_3/R vdd DFFSR_20/D gnd vdd DFFSR
XDFFSR_97 INVX4_9/A DFFSR_7/CLK DFFSR_99/R vdd DFFSR_97/D gnd vdd DFFSR
XCLKBUF1_51 CLKBUF1_3/A gnd DFFSR_6/CLK vdd CLKBUF1
XCLKBUF1_40 CLKBUF1_9/A gnd CLKBUF1_40/Y vdd CLKBUF1
XDFFSR_75 DFFSR_75/Q CLKBUF1_8/A DFFSR_2/R vdd DFFSR_75/D gnd vdd DFFSR
XDFFSR_86 DFFSR_86/Q DFFSR_86/CLK DFFSR_95/R vdd DFFSR_86/D gnd vdd DFFSR
XCLKBUF1_62 wb_clk_i gnd DFFSR_30/CLK vdd CLKBUF1
XINVX1_125 NOR3X1_6/B gnd INVX1_125/Y vdd INVX1
XINVX1_158 XOR2X1_3/B gnd INVX1_158/Y vdd INVX1
XINVX1_136 OR2X2_3/B gnd INVX1_136/Y vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XAOI21X1_118 MUX2X1_8/A OAI21X1_391/B BUFX4_264/Y gnd OAI21X1_391/C vdd AOI21X1
XAOI21X1_107 BUFX4_266/Y OAI21X1_378/Y BUFX4_249/Y gnd AOI22X1_48/D vdd AOI21X1
XAOI21X1_129 BUFX4_261/Y OAI21X1_402/Y BUFX4_245/Y gnd AOI22X1_57/D vdd AOI21X1
XFILL_23_0_1 gnd vdd FILL
XINVX4_11 INVX4_11/A gnd INVX4_11/Y vdd INVX4
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XDFFSR_109 INVX2_47/A CLKBUF1_5/Y vdd DFFSR_113/S DFFSR_109/D gnd vdd DFFSR
XBUFX4_264 BUFX4_268/A gnd BUFX4_264/Y vdd BUFX4
XBUFX4_231 INVX8_18/Y gnd BUFX4_231/Y vdd BUFX4
XBUFX4_220 BUFX4_220/A gnd BUFX4_220/Y vdd BUFX4
XBUFX4_275 BUFX4_277/A gnd MUX2X1_38/A vdd BUFX4
XBUFX4_253 BUFX4_255/A gnd BUFX4_253/Y vdd BUFX4
XBUFX4_242 BUFX4_242/A gnd INVX8_6/A vdd BUFX4
XNOR2X1_42 INVX1_70/Y AND2X2_5/Y gnd NOR2X1_42/Y vdd NOR2X1
XNAND3X1_42 INVX4_10/A OR2X2_3/B INVX4_9/A gnd OAI22X1_47/C vdd NAND3X1
XNOR2X1_31 INVX2_31/A INVX2_32/A gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_53 OR2X2_8/B INVX2_49/Y gnd INVX1_83/A vdd NOR2X1
XNOR2X1_64 INVX1_90/Y NOR2X1_64/B gnd NOR2X1_64/Y vdd NOR2X1
XNAND3X1_53 AND2X2_3/B OAI21X1_95/Y BUFX4_129/Y gnd OAI21X1_96/C vdd NAND3X1
XNOR2X1_20 NOR2X1_1/B INVX8_5/A gnd INVX8_15/A vdd NOR2X1
XNAND3X1_86 NAND3X1_86/A NAND3X1_86/B NAND3X1_86/C gnd DFFSR_95/D vdd NAND3X1
XNAND3X1_75 NAND3X1_75/A AOI22X1_8/Y AOI22X1_7/Y gnd DFFSR_84/D vdd NAND3X1
XNAND3X1_31 AND2X2_1/B OAI21X1_57/Y BUFX4_95/Y gnd OAI21X1_58/C vdd NAND3X1
XNAND3X1_97 BUFX4_64/Y NAND3X1_97/B NAND3X1_97/C gnd NAND3X1_97/Y vdd NAND3X1
XNAND3X1_64 AND2X2_1/B NAND3X1_64/B BUFX4_129/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_20 BUFX4_199/Y OAI21X1_35/Y BUFX4_96/Y gnd OAI21X1_36/C vdd NAND3X1
XNOR2X1_75 NOR2X1_75/A NOR2X1_75/B gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_86 INVX1_34/A NOR2X1_87/B gnd NOR2X1_86/Y vdd NOR2X1
XNOR2X1_97 INVX1_18/A NOR2X1_98/B gnd NOR2X1_97/Y vdd NOR2X1
XNAND2X1_8 BUFX4_86/Y wb_dat_i[31] gnd NAND2X1_8/Y vdd NAND2X1
XNOR2X1_176 INVX8_19/Y NOR2X1_193/B gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_165 OR2X2_13/B NOR2X1_189/B gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_110 INVX2_141/A NOR2X1_88/B gnd OAI22X1_66/C vdd NOR2X1
XNOR2X1_154 INVX2_158/Y INVX2_160/Y gnd NOR2X1_154/Y vdd NOR2X1
XNOR2X1_143 INVX1_48/A NOR2X1_79/B gnd OAI22X1_82/C vdd NOR2X1
XNOR2X1_132 INVX2_104/A NOR2X1_96/B gnd OAI22X1_77/C vdd NOR2X1
XNOR2X1_121 INVX2_77/A BUFX4_179/Y gnd OAI22X1_71/B vdd NOR2X1
XNOR2X1_198 INVX8_18/A NOR2X1_198/B gnd INVX1_154/A vdd NOR2X1
XOAI21X1_638 INVX1_113/Y BUFX4_25/Y OAI21X1_638/C gnd OAI21X1_638/Y vdd OAI21X1
XOAI21X1_649 BUFX4_121/Y INVX8_20/Y MUX2X1_38/Y gnd OAI21X1_650/C vdd OAI21X1
XOAI21X1_627 OAI21X1_627/A BUFX4_2/Y OAI21X1_627/C gnd DFFSR_132/D vdd OAI21X1
XOAI21X1_605 INVX1_105/Y BUFX4_187/Y OAI21X1_605/C gnd OAI21X1_605/Y vdd OAI21X1
XNOR2X1_187 BUFX4_251/Y INVX1_145/A gnd AND2X2_17/A vdd NOR2X1
XOAI21X1_616 OAI21X1_616/A BUFX4_7/Y OAI21X1_616/C gnd DFFSR_135/D vdd OAI21X1
XINVX1_78 OR2X2_2/A gnd INVX1_78/Y vdd INVX1
XINVX1_67 INVX2_35/A gnd INVX1_67/Y vdd INVX1
XINVX1_89 OR2X2_4/B gnd INVX1_89/Y vdd INVX1
XINVX1_45 INVX2_81/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_23 INVX2_94/A gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND3X1_272 INVX1_129/Y INVX2_151/A NAND3X1_272/C gnd NAND3X1_273/B vdd NAND3X1
XNAND3X1_261 OAI21X1_236/Y XNOR2X1_9/Y INVX1_131/A gnd AOI21X1_72/B vdd NAND3X1
XNAND3X1_250 BUFX4_64/Y NAND3X1_250/B NAND3X1_250/C gnd AOI21X1_58/B vdd NAND3X1
XFILL_22_6_0 gnd vdd FILL
XOAI22X1_18 INVX8_5/A INVX1_35/Y INVX8_2/A INVX2_28/Y gnd AOI21X1_6/C vdd OAI22X1
XOAI22X1_29 INVX8_1/A INVX2_3/Y INVX2_32/Y INVX8_4/A gnd NOR2X1_11/A vdd OAI22X1
XOAI21X1_424 BUFX4_231/Y OAI21X1_424/B BUFX4_43/Y gnd OAI22X1_85/D vdd OAI21X1
XOAI21X1_413 BUFX4_52/Y BUFX4_125/Y NOR2X1_147/Y gnd NOR2X1_189/B vdd OAI21X1
XOAI21X1_468 NOR2X1_174/Y INVX2_87/Y BUFX4_231/Y gnd OAI21X1_468/Y vdd OAI21X1
XOAI21X1_479 BUFX4_232/Y OAI21X1_479/B BUFX4_41/Y gnd OAI22X1_94/D vdd OAI21X1
XOAI21X1_435 INVX2_141/Y BUFX4_89/Y OAI21X1_525/C gnd OAI21X1_436/B vdd OAI21X1
XOAI21X1_446 BUFX4_158/Y OAI21X1_446/B OAI21X1_446/C gnd AOI22X1_63/C vdd OAI21X1
XOAI21X1_402 INVX2_64/Y MUX2X1_47/S OAI21X1_573/C gnd OAI21X1_402/Y vdd OAI21X1
XOAI21X1_457 BUFX4_53/Y BUFX4_126/Y NOR2X1_159/Y gnd INVX1_147/A vdd OAI21X1
XFILL_5_7_0 gnd vdd FILL
XFILL_13_6_0 gnd vdd FILL
XOAI21X1_84 AND2X2_2/Y INVX2_26/Y OAI21X1_84/C gnd DFFSR_36/D vdd OAI21X1
XOAI21X1_73 BUFX4_29/Y BUFX4_23/Y OAI21X1_73/C gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_51 INVX2_11/Y BUFX4_108/Y OAI21X1_79/C gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_95 INVX2_32/Y BUFX4_26/Y OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_62 BUFX4_101/Y INVX2_16/Y OAI21X1_62/C gnd DFFSR_7/D vdd OAI21X1
XOAI21X1_40 OAI21X1_2/A INVX2_5/Y OAI21X1_40/C gnd DFFSR_12/D vdd OAI21X1
XOAI21X1_210 XNOR2X1_7/Y BUFX4_181/Y NAND2X1_95/Y gnd BUFX4_207/A vdd OAI21X1
XOAI21X1_221 AND2X2_11/Y NOR2X1_65/Y INVX2_55/Y gnd AOI21X1_41/B vdd OAI21X1
XOAI21X1_243 XNOR2X1_12/B XNOR2X1_11/Y NOR2X1_70/Y gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_232 INVX1_82/Y NOR2X1_52/Y OAI21X1_232/C gnd DFFSR_244/D vdd OAI21X1
XAND2X2_10 OR2X2_4/A AND2X2_10/B gnd AND2X2_10/Y vdd AND2X2
XOAI21X1_254 INVX1_127/Y INVX4_8/Y OAI21X1_254/C gnd OAI21X1_254/Y vdd OAI21X1
XOAI21X1_276 NOR2X1_82/B INVX1_100/A BUFX4_38/Y gnd OAI22X1_58/A vdd OAI21X1
XAND2X2_21 MUX2X1_34/A AND2X2_21/B gnd AND2X2_21/Y vdd AND2X2
XOAI21X1_287 INVX1_56/A NOR2X1_84/B BUFX4_168/Y gnd OAI22X1_61/A vdd OAI21X1
XOAI21X1_265 INVX2_86/A NOR2X1_84/B BUFX4_77/Y gnd OAI22X1_53/D vdd OAI21X1
XOAI21X1_298 INVX2_139/A NOR2X1_88/B BUFX4_77/Y gnd OAI22X1_65/D vdd OAI21X1
XNAND2X1_260 INVX4_9/A AND2X2_10/Y gnd OAI21X1_707/C vdd NAND2X1
XDFFSR_76 DFFSR_76/Q DFFSR_1/CLK DFFSR_93/R vdd DFFSR_76/D gnd vdd DFFSR
XDFFSR_98 MUX2X1_1/A DFFSR_98/CLK DFFSR_99/R vdd DFFSR_98/D gnd vdd DFFSR
XDFFSR_65 DFFSR_65/Q CLKBUF1_2/Y DFFSR_93/R vdd DFFSR_65/D gnd vdd DFFSR
XDFFSR_54 INVX2_46/A DFFSR_99/CLK DFFSR_93/R vdd DFFSR_54/D gnd vdd DFFSR
XDFFSR_43 MUX2X1_1/S DFFSR_58/CLK DFFSR_80/R vdd DFFSR_43/D gnd vdd DFFSR
XDFFSR_87 DFFSR_87/Q DFFSR_87/CLK DFFSR_96/R vdd DFFSR_87/D gnd vdd DFFSR
XDFFSR_21 INVX1_13/A DFFSR_96/CLK DFFSR_96/R vdd DFFSR_21/D gnd vdd DFFSR
XDFFSR_32 INVX1_8/A DFFSR_92/CLK DFFSR_3/R vdd DFFSR_32/D gnd vdd DFFSR
XDFFSR_10 INVX2_3/A DFFSR_85/CLK DFFSR_9/R vdd DFFSR_10/D gnd vdd DFFSR
XCLKBUF1_41 CLKBUF1_61/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XCLKBUF1_30 CLKBUF1_64/Y gnd DFFSR_41/CLK vdd CLKBUF1
XCLKBUF1_63 wb_clk_i gnd CLKBUF1_63/Y vdd CLKBUF1
XCLKBUF1_52 CLKBUF1_63/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XFILL_27_5_0 gnd vdd FILL
XFILL_2_5_0 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_126 INVX1_126/A gnd NOR3X1_6/C vdd INVX1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_115 MUX2X1_41/B gnd MUX2X1_42/B vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XFILL_18_5_0 gnd vdd FILL
XAOI21X1_119 BUFX4_263/Y OAI21X1_392/Y BUFX4_243/Y gnd AOI22X1_52/D vdd AOI21X1
XAOI21X1_108 INVX2_106/Y INVX1_141/Y BUFX4_268/Y gnd AOI21X1_109/A vdd AOI21X1
XINVX4_12 INVX4_12/A gnd INVX4_12/Y vdd INVX4
XBUFX4_276 BUFX4_277/A gnd MUX2X1_34/A vdd BUFX4
XBUFX4_210 INVX8_8/Y gnd DFFSR_80/R vdd BUFX4
XBUFX4_243 BUFX4_250/A gnd BUFX4_243/Y vdd BUFX4
XBUFX4_232 INVX8_18/Y gnd BUFX4_232/Y vdd BUFX4
XBUFX4_254 BUFX4_255/A gnd BUFX4_254/Y vdd BUFX4
XBUFX4_221 BUFX4_228/A gnd NOR2X1_98/B vdd BUFX4
XBUFX4_265 BUFX4_268/A gnd BUFX4_265/Y vdd BUFX4
XFILL_24_3_0 gnd vdd FILL
XNAND3X1_21 BUFX4_202/Y OAI21X1_37/Y BUFX4_97/Y gnd OAI21X1_38/C vdd NAND3X1
XNAND3X1_32 BUFX4_200/Y OAI21X1_59/Y BUFX4_97/Y gnd OAI21X1_60/C vdd NAND3X1
XNAND3X1_10 AND2X2_1/B OAI21X1_15/Y BUFX4_98/Y gnd OAI21X1_16/C vdd NAND3X1
XFILL_7_4_0 gnd vdd FILL
XNOR2X1_43 INVX1_72/Y NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_76 NOR2X1_76/A NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_54 NOR2X1_54/A AND2X2_8/Y gnd INVX1_84/A vdd NOR2X1
XNOR2X1_32 INVX2_37/A INVX2_36/A gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_21 INVX2_47/A INVX1_74/A gnd INVX1_75/A vdd NOR2X1
XNAND3X1_54 AND2X2_2/B OAI21X1_97/Y BUFX4_131/Y gnd OAI21X1_98/C vdd NAND3X1
XNOR2X1_65 MUX2X1_6/Y BUFX4_66/Y gnd NOR2X1_65/Y vdd NOR2X1
XNAND3X1_65 BUFX4_200/Y NAND3X1_65/B BUFX4_130/Y gnd NAND3X1_65/Y vdd NAND3X1
XNAND3X1_43 OAI21X1_77/Y NAND3X1_7/A INVX8_2/Y gnd OAI21X1_78/C vdd NAND3X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_87 INVX2_98/A NOR2X1_87/B gnd NOR2X1_87/Y vdd NOR2X1
XNAND3X1_76 NAND3X1_76/A NAND3X1_76/B AOI22X1_9/Y gnd DFFSR_85/D vdd NAND3X1
XNAND3X1_87 NAND3X1_87/A NAND3X1_87/B NAND3X1_87/C gnd DFFSR_96/D vdd NAND3X1
XNAND3X1_98 INVX1_95/Y BUFX4_50/Y BUFX4_137/Y gnd NAND3X1_98/Y vdd NAND3X1
XFILL_15_3_0 gnd vdd FILL
XNOR2X1_98 NOR2X1_98/A NOR2X1_98/B gnd NOR2X1_98/Y vdd NOR2X1
XNAND2X1_9 wb_dat_i[16] NAND2X1_9/B gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_166 OR2X2_13/B NOR2X1_191/B gnd NOR2X1_166/Y vdd NOR2X1
XNOR2X1_100 INVX2_132/A NOR2X1_99/B gnd OAI22X1_61/C vdd NOR2X1
XNOR2X1_111 XOR2X1_6/Y NOR2X1_94/B gnd INVX2_159/A vdd NOR2X1
XNOR2X1_144 XOR2X1_6/Y NOR2X1_74/B gnd INVX2_157/A vdd NOR2X1
XNOR2X1_199 INVX4_11/Y INVX1_154/Y gnd NOR2X1_199/Y vdd NOR2X1
XNOR2X1_177 INVX8_19/Y NOR2X1_195/B gnd NOR2X1_177/Y vdd NOR2X1
XNOR2X1_188 BUFX4_127/Y INVX8_22/Y gnd BUFX4_260/A vdd NOR2X1
XNOR2X1_133 INVX1_60/A NOR2X1_78/B gnd OAI22X1_77/B vdd NOR2X1
XNOR2X1_122 INVX2_75/A NOR2X1_71/A gnd OAI22X1_72/B vdd NOR2X1
XNOR2X1_155 INVX2_159/Y INVX2_160/Y gnd NOR2X1_155/Y vdd NOR2X1
XOAI21X1_639 AND2X2_27/B INVX1_113/A BUFX4_166/Y gnd OAI21X1_640/B vdd OAI21X1
XOAI21X1_628 BUFX4_121/Y INVX8_20/Y MUX2X1_32/Y gnd OAI21X1_629/C vdd OAI21X1
XOAI21X1_617 INVX1_114/Y BUFX4_190/Y OAI21X1_617/C gnd OAI21X1_617/Y vdd OAI21X1
XOAI21X1_606 BUFX4_127/Y INVX8_22/Y AND2X2_19/A gnd NOR2X1_238/B vdd OAI21X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_46 INVX2_79/A gnd INVX1_46/Y vdd INVX1
XINVX1_57 INVX2_87/A gnd INVX1_57/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XNAND3X1_273 BUFX4_272/Y NAND3X1_273/B OAI21X1_260/Y gnd AOI21X1_77/B vdd NAND3X1
XFILL_30_1_0 gnd vdd FILL
XNAND3X1_262 INVX2_48/A OR2X2_4/B NOR3X1_5/Y gnd INVX1_126/A vdd NAND3X1
XNAND3X1_251 INVX1_107/Y NAND3X1_251/B OAI21X1_231/Y gnd NAND3X1_252/C vdd NAND3X1
XNAND3X1_240 INVX2_146/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_241/C vdd NAND3X1
XFILL_22_6_1 gnd vdd FILL
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 NOR2X1_165/Y INVX2_88/Y BUFX4_231/Y gnd OAI21X1_414/Y vdd OAI21X1
XOAI21X1_403 BUFX4_155/Y OAI21X1_403/B OAI21X1_403/C gnd AOI22X1_58/C vdd OAI21X1
XOAI22X1_19 OAI22X1_7/A INVX1_37/Y INVX1_36/Y OAI22X1_7/D gnd NOR2X1_8/B vdd OAI22X1
XOAI21X1_469 INVX2_87/Y BUFX4_24/Y OAI21X1_630/C gnd OAI21X1_470/B vdd OAI21X1
XOAI21X1_436 BUFX4_232/Y OAI21X1_436/B BUFX4_41/Y gnd OAI22X1_88/D vdd OAI21X1
XOAI21X1_425 BUFX4_55/Y BUFX4_125/Y INVX1_142/A gnd NOR2X1_195/B vdd OAI21X1
XOAI21X1_447 INVX2_138/Y BUFX4_188/Y OAI21X1_609/C gnd OAI21X1_448/B vdd OAI21X1
XOAI21X1_458 BUFX4_158/Y OAI21X1_458/B OAI21X1_458/C gnd AOI22X1_65/C vdd OAI21X1
XFILL_5_7_1 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_41 INVX2_6/Y BUFX4_20/Y OAI21X1_71/C gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_52 OAI21X1_8/A INVX2_11/Y OAI21X1_52/C gnd DFFSR_2/D vdd OAI21X1
XOAI21X1_63 INVX2_17/Y MUX2X1_47/S OAI21X1_91/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_30 BUFX4_102/Y INVX1_15/Y OAI21X1_30/C gnd DFFSR_23/D vdd OAI21X1
XOAI21X1_74 AND2X2_2/Y BUFX4_29/Y OAI21X1_74/C gnd DFFSR_46/D vdd OAI21X1
XOAI21X1_96 AND2X2_3/Y INVX2_32/Y OAI21X1_96/C gnd DFFSR_56/D vdd OAI21X1
XOAI21X1_85 INVX2_27/Y MUX2X1_35/S OAI21X1_85/C gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_244 OAI21X1_244/A OAI21X1_244/B AOI21X1_69/Y gnd NOR2X1_76/B vdd OAI21X1
XOAI21X1_233 OR2X2_7/A OR2X2_7/B INVX4_7/Y gnd AOI21X1_61/A vdd OAI21X1
XOAI21X1_211 NOR2X1_49/B INVX4_7/A INVX2_48/A gnd AND2X2_10/B vdd OAI21X1
XOAI21X1_255 AOI21X1_66/Y INVX1_128/A OR2X2_9/B gnd OAI21X1_256/A vdd OAI21X1
XOAI21X1_200 BUFX2_80/A NOR2X1_256/B OAI21X1_200/C gnd NOR3X1_4/B vdd OAI21X1
XOAI21X1_222 NOR2X1_67/Y NOR2X1_66/Y INVX2_55/A gnd AOI21X1_41/A vdd OAI21X1
XAND2X2_11 BUFX4_66/Y AND2X2_11/B gnd AND2X2_11/Y vdd AND2X2
XOAI21X1_277 NOR2X1_99/B MUX2X1_25/B BUFX4_33/Y gnd OAI22X1_58/D vdd OAI21X1
XOAI21X1_288 INVX2_128/A NOR2X1_84/B BUFX4_77/Y gnd OAI22X1_61/D vdd OAI21X1
XOAI21X1_266 NOR2X1_82/B INVX1_101/A BUFX4_38/Y gnd OAI22X1_54/A vdd OAI21X1
XOAI21X1_299 NOR2X1_87/B INVX1_121/A BUFX4_37/Y gnd OAI22X1_66/A vdd OAI21X1
XAND2X2_22 MUX2X1_42/A AND2X2_22/B gnd AND2X2_22/Y vdd AND2X2
XNAND2X1_261 INVX2_52/A INVX4_10/Y gnd OAI21X1_708/C vdd NAND2X1
XNAND2X1_250 INVX4_12/A NOR2X1_246/Y gnd OAI21X1_686/B vdd NAND2X1
XDFFSR_99 OR2X2_1/B DFFSR_99/CLK DFFSR_99/R vdd DFFSR_99/D gnd vdd DFFSR
XDFFSR_66 DFFSR_66/Q DFFSR_6/CLK DFFSR_93/R vdd DFFSR_66/D gnd vdd DFFSR
XDFFSR_44 DFFSR_44/Q CLKBUF1_3/A DFFSR_80/R vdd DFFSR_44/D gnd vdd DFFSR
XDFFSR_55 INVX2_31/A DFFSR_55/CLK DFFSR_63/R vdd DFFSR_55/D gnd vdd DFFSR
XDFFSR_33 OR2X2_8/B DFFSR_93/CLK DFFSR_80/R vdd DFFSR_33/D gnd vdd DFFSR
XDFFSR_77 DFFSR_77/Q DFFSR_2/CLK DFFSR_2/R vdd DFFSR_77/D gnd vdd DFFSR
XDFFSR_11 INVX2_4/A DFFSR_71/CLK DFFSR_7/R vdd DFFSR_11/D gnd vdd DFFSR
XDFFSR_22 INVX1_14/A DFFSR_82/CLK DFFSR_95/R vdd DFFSR_22/D gnd vdd DFFSR
XDFFSR_88 DFFSR_88/Q DFFSR_88/CLK DFFSR_95/R vdd DFFSR_88/D gnd vdd DFFSR
XCLKBUF1_64 wb_clk_i gnd CLKBUF1_64/Y vdd CLKBUF1
XCLKBUF1_53 wb_clk_i gnd CLKBUF1_7/A vdd CLKBUF1
XCLKBUF1_20 CLKBUF1_63/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_42 DFFSR_30/CLK gnd DFFSR_83/CLK vdd CLKBUF1
XCLKBUF1_31 CLKBUF1_6/A gnd DFFSR_86/CLK vdd CLKBUF1
XFILL_27_5_1 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_116 MUX2X1_33/B gnd MUX2X1_34/B vdd INVX1
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XFILL_10_4_1 gnd vdd FILL
XINVX1_127 OR2X2_5/B gnd INVX1_127/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XINVX1_149 BUFX4_36/Y gnd INVX1_149/Y vdd INVX1
XFILL_18_5_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 AOI21X1_109/A NAND2X1_178/Y AND2X2_15/Y gnd OAI21X1_381/A vdd AOI21X1
XBUFX4_200 NOR2X1_1/Y gnd BUFX4_200/Y vdd BUFX4
XBUFX4_211 INVX8_8/Y gnd DFFSR_95/R vdd BUFX4
XBUFX4_233 INVX8_18/Y gnd BUFX4_233/Y vdd BUFX4
XBUFX4_244 BUFX4_250/A gnd BUFX4_244/Y vdd BUFX4
XBUFX4_266 BUFX4_268/A gnd BUFX4_266/Y vdd BUFX4
XBUFX4_255 BUFX4_255/A gnd BUFX4_255/Y vdd BUFX4
XBUFX4_277 BUFX4_277/A gnd MUX2X1_42/A vdd BUFX4
XBUFX4_222 BUFX4_228/A gnd BUFX4_222/Y vdd BUFX4
XFILL_24_3_1 gnd vdd FILL
XNAND3X1_55 BUFX4_202/Y OAI21X1_99/Y BUFX4_131/Y gnd NAND3X1_55/Y vdd NAND3X1
XNAND3X1_66 BUFX4_202/Y NAND3X1_66/B AND2X2_3/A gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_44 OAI21X1_79/Y NAND3X1_7/A INVX8_2/Y gnd OAI21X1_80/C vdd NAND3X1
XNAND3X1_33 AND2X2_3/B OAI21X1_61/Y BUFX4_97/Y gnd OAI21X1_62/C vdd NAND3X1
XNAND3X1_11 NAND3X1_9/A OAI21X1_17/Y BUFX4_94/Y gnd OAI21X1_18/C vdd NAND3X1
XFILL_7_4_1 gnd vdd FILL
XNAND3X1_22 BUFX4_199/Y OAI21X1_39/Y BUFX4_96/Y gnd OAI21X1_40/C vdd NAND3X1
XNAND3X1_88 XOR2X1_1/A INVX1_65/Y AND2X2_5/A gnd NOR2X1_29/B vdd NAND3X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_22 NOR3X1_2/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_44 NOR3X1_2/B NOR3X1_3/C gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_11 NOR2X1_11/A NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_55 XNOR2X1_3/Y INVX1_83/Y gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_66 MUX2X1_7/Y NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_99 INVX1_55/A NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_88 INVX1_33/A NOR2X1_88/B gnd NOR2X1_88/Y vdd NOR2X1
XNOR2X1_77 INVX2_95/A NOR2X1_87/B gnd NOR2X1_77/Y vdd NOR2X1
XNAND3X1_77 NAND3X1_77/A NAND3X1_77/B NAND3X1_77/C gnd DFFSR_86/D vdd NAND3X1
XNAND3X1_99 INVX2_63/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_99/Y vdd NAND3X1
XFILL_30_1 gnd vdd FILL
XNOR2X1_178 INVX8_19/Y NOR2X1_196/B gnd NOR2X1_178/Y vdd NOR2X1
XNOR2X1_101 INVX1_54/A NOR2X1_93/B gnd OAI22X1_62/B vdd NOR2X1
XNOR2X1_167 OR2X2_13/B NOR2X1_193/B gnd NOR2X1_167/Y vdd NOR2X1
XNOR2X1_189 INVX8_18/A NOR2X1_189/B gnd INVX1_150/A vdd NOR2X1
XNOR2X1_145 BUFX4_125/Y BUFX4_55/Y gnd BUFX4_268/A vdd NOR2X1
XNOR2X1_134 INVX2_105/A BUFX4_222/Y gnd OAI22X1_78/B vdd NOR2X1
XNOR2X1_112 INVX2_61/A NOR2X1_78/B gnd OAI22X1_67/C vdd NOR2X1
XNOR2X1_123 INVX2_78/A NOR2X1_71/A gnd OAI22X1_72/C vdd NOR2X1
XMUX2X1_40 MUX2X1_48/A INVX1_95/Y MUX2X1_40/S gnd MUX2X1_40/Y vdd MUX2X1
XNOR2X1_156 NOR2X1_75/A INVX2_154/A gnd NOR2X1_156/Y vdd NOR2X1
XOAI21X1_629 BUFX4_163/Y MUX2X1_31/Y OAI21X1_629/C gnd DFFSR_130/D vdd OAI21X1
XOAI21X1_607 AND2X2_22/B INVX1_105/A BUFX4_161/Y gnd OAI21X1_608/B vdd OAI21X1
XOAI21X1_618 BUFX4_127/Y INVX8_22/Y NOR2X1_203/Y gnd NOR2X1_241/B vdd OAI21X1
XINVX1_47 INVX2_83/A gnd INVX1_47/Y vdd INVX1
XINVX1_58 INVX2_89/A gnd INVX1_58/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_69 INVX2_43/A gnd INVX1_69/Y vdd INVX1
XNAND3X1_230 MUX2X1_28/B BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_232/B vdd NAND3X1
XNAND3X1_241 BUFX4_204/Y NAND3X1_241/B NAND3X1_241/C gnd AOI21X1_57/A vdd NAND3X1
XFILL_30_1_1 gnd vdd FILL
XNAND3X1_263 INVX2_52/A NAND3X1_263/B OAI21X1_238/Y gnd INVX2_151/A vdd NAND3X1
XNAND3X1_252 NOR2X1_52/Y NAND3X1_252/B NAND3X1_252/C gnd OAI21X1_232/C vdd NAND3X1
XNAND3X1_274 OR2X2_10/A OAI21X1_279/Y OAI21X1_302/Y gnd OAI21X1_345/A vdd NAND3X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_415 INVX2_88/Y BUFX4_91/Y OAI21X1_511/C gnd OAI21X1_416/B vdd OAI21X1
XOAI21X1_426 NOR2X1_168/Y INVX2_117/Y BUFX4_233/Y gnd OAI21X1_426/Y vdd OAI21X1
XOAI21X1_448 BUFX4_143/Y OAI21X1_448/B BUFX4_249/Y gnd AOI22X1_63/D vdd OAI21X1
XOAI21X1_404 INVX2_124/Y BUFX4_106/Y OAI21X1_575/C gnd OAI21X1_404/Y vdd OAI21X1
XOAI21X1_437 BUFX4_53/Y BUFX4_126/Y NOR2X1_153/Y gnd OR2X2_11/A vdd OAI21X1
XDFFSR_250 INVX2_48/A DFFSR_70/CLK BUFX4_15/Y vdd DFFSR_250/D gnd vdd DFFSR
XOAI21X1_459 INVX2_91/Y NAND2X1_9/B OAI21X1_621/C gnd OAI21X1_460/B vdd OAI21X1
XFILL_29_2_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XINVX2_90 INVX2_90/A gnd INVX2_90/Y vdd INVX2
XOAI21X1_75 INVX1_17/Y BUFX4_24/Y OAI21X1_93/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_42 OAI21X1_8/A INVX2_6/Y OAI21X1_42/C gnd DFFSR_13/D vdd OAI21X1
XOAI21X1_86 AND2X2_2/Y INVX2_27/Y OAI21X1_86/C gnd DFFSR_37/D vdd OAI21X1
XOAI21X1_64 BUFX4_101/Y INVX2_17/Y OAI21X1_64/C gnd DFFSR_8/D vdd OAI21X1
XOAI21X1_31 INVX1_16/Y BUFX4_185/Y OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_20 BUFX4_102/Y INVX1_10/Y OAI21X1_20/C gnd DFFSR_18/D vdd OAI21X1
XOAI21X1_53 INVX2_12/Y MUX2X1_37/S OAI21X1_81/C gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_97 INVX2_33/Y BUFX4_19/Y OAI21X1_97/C gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_201 INVX4_2/A INVX4_4/Y INVX1_87/A gnd XNOR2X1_5/A vdd OAI21X1
XOAI21X1_256 OAI21X1_256/A NOR2X1_76/Y OAI21X1_256/C gnd BUFX4_179/A vdd OAI21X1
XOAI21X1_234 OAI21X1_235/A INVX4_8/Y INVX4_2/A gnd OAI21X1_235/C vdd OAI21X1
XOAI21X1_245 INVX1_89/Y INVX4_8/Y NOR2X1_73/B gnd AOI21X1_71/C vdd OAI21X1
XOAI21X1_289 NOR2X1_82/B MUX2X1_33/B BUFX4_38/Y gnd OAI22X1_62/A vdd OAI21X1
XOAI21X1_278 OAI22X1_57/Y OAI22X1_58/Y INVX2_155/Y gnd OAI21X1_278/Y vdd OAI21X1
XOAI21X1_223 AOI21X1_41/Y NOR3X1_4/Y INVX4_5/Y gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_267 NOR2X1_82/B MUX2X1_19/B BUFX4_33/Y gnd OAI22X1_54/D vdd OAI21X1
XOAI21X1_212 XOR2X1_4/Y BUFX4_180/Y NAND2X1_96/Y gnd BUFX4_85/A vdd OAI21X1
XAND2X2_12 INVX2_151/A AND2X2_12/B gnd AND2X2_12/Y vdd AND2X2
XAND2X2_23 INVX8_14/A AND2X2_23/B gnd AND2X2_23/Y vdd AND2X2
XNAND2X1_262 NOR2X1_51/A INVX4_10/A gnd OAI21X1_711/B vdd NAND2X1
XNAND2X1_240 BUFX4_3/Y OAI21X1_651/Y gnd OAI21X1_653/C vdd NAND2X1
XNAND2X1_251 INVX4_11/A NOR2X1_250/Y gnd OAI21X1_688/B vdd NAND2X1
XDFFSR_12 INVX2_5/A DFFSR_87/CLK DFFSR_96/R vdd DFFSR_12/D gnd vdd DFFSR
XDFFSR_45 INVX2_22/A CLKBUF1_3/A DFFSR_80/R vdd DFFSR_45/D gnd vdd DFFSR
XDFFSR_34 INVX4_3/A CLKBUF1_5/Y DFFSR_80/R vdd DFFSR_34/D gnd vdd DFFSR
XDFFSR_78 DFFSR_78/Q CLKBUF1_9/Y DFFSR_2/R vdd DFFSR_78/D gnd vdd DFFSR
XDFFSR_56 INVX2_32/A DFFSR_71/CLK DFFSR_7/R vdd DFFSR_56/D gnd vdd DFFSR
XDFFSR_23 INVX1_15/A DFFSR_83/CLK DFFSR_95/R vdd DFFSR_23/D gnd vdd DFFSR
XDFFSR_67 DFFSR_67/Q DFFSR_82/CLK DFFSR_96/R vdd DFFSR_67/D gnd vdd DFFSR
XDFFSR_89 DFFSR_89/Q CLKBUF1_4/A DFFSR_3/R vdd DFFSR_89/D gnd vdd DFFSR
XCLKBUF1_54 wb_clk_i gnd CLKBUF1_54/Y vdd CLKBUF1
XCLKBUF1_43 CLKBUF1_3/A gnd DFFSR_8/CLK vdd CLKBUF1
XCLKBUF1_65 wb_clk_i gnd CLKBUF1_9/A vdd CLKBUF1
XCLKBUF1_21 CLKBUF1_9/A gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_10 CLKBUF1_7/A gnd CLKBUF1_10/Y vdd CLKBUF1
XCLKBUF1_32 CLKBUF1_4/A gnd DFFSR_71/CLK vdd CLKBUF1
XFILL_26_0_1 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XINVX1_128 INVX1_128/A gnd NOR2X1_76/A vdd INVX1
XINVX1_117 MUX2X1_21/B gnd MUX2X1_22/B vdd INVX1
XINVX1_106 MUX2X1_37/B gnd MUX2X1_38/B vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_20_7_0 gnd vdd FILL
XFILL_11_7_0 gnd vdd FILL
XBUFX4_212 INVX8_8/Y gnd DFFSR_93/R vdd BUFX4
XBUFX4_234 INVX8_18/Y gnd BUFX4_234/Y vdd BUFX4
XBUFX4_201 NOR2X1_1/Y gnd AND2X2_3/B vdd BUFX4
XBUFX4_245 BUFX4_250/A gnd BUFX4_245/Y vdd BUFX4
XBUFX4_223 BUFX4_228/A gnd NOR2X1_71/A vdd BUFX4
XBUFX4_267 BUFX4_268/A gnd BUFX4_267/Y vdd BUFX4
XBUFX4_256 BUFX4_260/A gnd INVX8_23/A vdd BUFX4
XNAND3X1_89 NOR2X1_30/Y NOR2X1_31/Y NOR2X1_32/Y gnd NOR2X1_33/B vdd NAND3X1
XNAND3X1_56 BUFX4_202/Y NAND3X1_56/B BUFX4_131/Y gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_23 BUFX4_200/Y OAI21X1_41/Y BUFX4_97/Y gnd OAI21X1_42/C vdd NAND3X1
XNAND3X1_67 BUFX4_202/Y NAND3X1_67/B AND2X2_3/A gnd NAND3X1_67/Y vdd NAND3X1
XNAND3X1_45 OAI21X1_81/Y NAND3X1_7/A INVX8_2/Y gnd OAI21X1_82/C vdd NAND3X1
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XNAND3X1_34 BUFX4_199/Y OAI21X1_63/Y BUFX4_96/Y gnd OAI21X1_64/C vdd NAND3X1
XNAND3X1_78 NAND3X1_78/A NAND3X1_78/B NAND3X1_78/C gnd DFFSR_87/D vdd NAND3X1
XNAND3X1_12 NAND3X1_9/A OAI21X1_19/Y BUFX4_93/Y gnd OAI21X1_20/C vdd NAND3X1
XNOR2X1_23 NOR3X1_3/A NOR2X1_23/B gnd INVX1_80/A vdd NOR2X1
XNOR2X1_45 OR2X2_2/A NOR3X1_3/C gnd NOR2X1_46/A vdd NOR2X1
XNOR2X1_34 INVX2_41/A INVX2_42/A gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_56 XNOR2X1_4/Y NOR2X1_56/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 MUX2X1_8/Y BUFX4_66/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_78 INVX2_93/A NOR2X1_78/B gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_89 INVX2_99/A NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_102 INVX2_130/A NOR2X1_93/B gnd OAI22X1_62/C vdd NOR2X1
XNOR2X1_124 INVX2_54/A NOR2X1_99/B gnd OAI22X1_73/C vdd NOR2X1
XMUX2X1_30 MUX2X1_42/A MUX2X1_30/B MUX2X1_30/S gnd MUX2X1_30/Y vdd MUX2X1
XMUX2X1_41 wb_dat_i[2] MUX2X1_41/B MUX2X1_41/S gnd MUX2X1_41/Y vdd MUX2X1
XNOR2X1_113 INVX2_65/A NOR2X1_78/B gnd OAI22X1_67/B vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XNOR2X1_179 INVX8_19/Y NOR2X1_198/B gnd NOR2X1_179/Y vdd NOR2X1
XNOR2X1_146 INVX2_157/Y NOR2X1_75/B gnd INVX1_140/A vdd NOR2X1
XNOR2X1_168 OR2X2_13/B NOR2X1_195/B gnd NOR2X1_168/Y vdd NOR2X1
XOAI21X1_619 AND2X2_24/B INVX1_114/A BUFX4_165/Y gnd OAI21X1_620/B vdd OAI21X1
XOAI21X1_608 AND2X2_22/Y OAI21X1_608/B OAI21X1_608/C gnd DFFSR_137/D vdd OAI21X1
XNOR2X1_135 INVX1_61/A NOR2X1_89/B gnd OAI22X1_78/C vdd NOR2X1
XNOR2X1_157 INVX2_157/Y INVX2_154/A gnd NOR2X1_157/Y vdd NOR2X1
XINVX1_59 INVX2_85/A gnd INVX1_59/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XFILL_25_6_0 gnd vdd FILL
XFILL_0_6_0 gnd vdd FILL
XFILL_8_7_0 gnd vdd FILL
XNAND3X1_264 INVX2_52/Y NAND3X1_264/B OAI21X1_239/Y gnd AND2X2_12/B vdd NAND3X1
XNAND3X1_275 INVX1_158/Y INVX4_6/Y NOR2X1_260/Y gnd NOR2X1_261/B vdd NAND3X1
XNAND3X1_253 OR2X2_5/A OR2X2_5/B INVX4_8/A gnd OR2X2_7/A vdd NAND3X1
XNAND3X1_231 INVX2_141/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_232/C vdd NAND3X1
XFILL_16_6_0 gnd vdd FILL
XNAND3X1_242 INVX1_122/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_244/B vdd NAND3X1
XNAND3X1_220 BUFX4_62/Y NAND3X1_220/B NAND3X1_220/C gnd AOI21X1_52/B vdd NAND3X1
XOAI21X1_416 BUFX4_231/Y OAI21X1_416/B BUFX4_43/Y gnd OAI22X1_83/D vdd OAI21X1
XOAI21X1_405 BUFX4_160/Y OAI21X1_405/B OAI21X1_405/C gnd AOI22X1_59/C vdd OAI21X1
XOAI21X1_427 INVX2_117/Y BUFX4_87/Y OAI21X1_520/C gnd OAI21X1_428/B vdd OAI21X1
XOAI21X1_438 BUFX4_157/Y OR2X2_11/Y OAI21X1_438/C gnd AOI22X1_62/C vdd OAI21X1
XOAI21X1_449 BUFX4_53/Y BUFX4_126/Y NOR2X1_156/Y gnd NOR2X1_202/B vdd OAI21X1
XDFFSR_251 OR2X2_4/B CLKBUF1_29/Y BUFX4_15/Y vdd DFFSR_251/D gnd vdd DFFSR
XDFFSR_240 INVX2_128/A CLKBUF1_60/Y BUFX4_8/Y vdd DFFSR_240/D gnd vdd DFFSR
XINVX2_80 INVX2_80/A gnd MUX2X1_6/B vdd INVX2
XINVX2_91 INVX2_91/A gnd INVX2_91/Y vdd INVX2
XOAI21X1_76 AND2X2_2/Y OAI21X1_76/B OAI21X1_76/C gnd DFFSR_41/D vdd OAI21X1
XOAI21X1_65 INVX2_18/Y BUFX4_19/Y OAI21X1_95/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_98 AND2X2_3/Y INVX2_33/Y OAI21X1_98/C gnd DFFSR_57/D vdd OAI21X1
XOAI21X1_10 OAI21X1_8/A INVX1_5/Y NAND3X1_7/Y gnd DFFSR_29/D vdd OAI21X1
XOAI21X1_87 INVX2_28/Y MUX2X1_37/S OAI21X1_87/C gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_43 INVX2_7/Y BUFX4_22/Y OAI21X1_73/C gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_32 BUFX4_102/Y INVX1_16/Y OAI21X1_32/C gnd DFFSR_24/D vdd OAI21X1
XOAI21X1_21 INVX1_11/Y BUFX4_189/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_54 OAI21X1_2/A INVX2_12/Y OAI21X1_54/C gnd DFFSR_3/D vdd OAI21X1
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_246 AOI21X1_72/Y INVX2_151/Y INVX1_129/Y gnd AOI21X1_73/B vdd OAI21X1
XOAI21X1_202 OR2X2_5/Y INVX4_2/A INVX4_7/A gnd AND2X2_9/B vdd OAI21X1
XOAI21X1_235 OAI21X1_235/A OAI21X1_251/C OAI21X1_235/C gnd XNOR2X1_9/A vdd OAI21X1
XAND2X2_13 AND2X2_13/A OR2X2_9/Y gnd NOR3X1_8/A vdd AND2X2
XOAI21X1_257 OR2X2_9/B OR2X2_9/A AND2X2_13/A gnd NOR3X1_9/B vdd OAI21X1
XOAI21X1_213 XOR2X1_5/Y BUFX4_181/Y NAND2X1_98/Y gnd BUFX4_66/A vdd OAI21X1
XOAI21X1_268 OAI22X1_53/Y OAI22X1_54/Y NOR2X1_72/Y gnd OAI21X1_268/Y vdd OAI21X1
XOAI21X1_279 OAI21X1_279/A OAI21X1_279/B NOR2X1_94/Y gnd OAI21X1_279/Y vdd OAI21X1
XOAI21X1_224 AOI21X1_44/Y AOI21X1_45/Y INVX4_5/Y gnd OAI21X1_224/Y vdd OAI21X1
XAND2X2_24 MUX2X1_42/A AND2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XNAND2X1_230 BUFX4_2/Y OAI21X1_617/Y gnd OAI21X1_620/C vdd NAND2X1
XNAND2X1_241 NOR2X1_239/Y INVX8_14/A gnd OAI21X1_652/C vdd NAND2X1
XNAND2X1_252 INVX4_12/A NOR2X1_250/Y gnd OAI21X1_690/B vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XFILL_13_4_0 gnd vdd FILL
XDFFSR_35 INVX4_4/A CLKBUF1_3/Y DFFSR_80/R vdd DFFSR_35/D gnd vdd DFFSR
XDFFSR_13 INVX2_6/A DFFSR_58/CLK DFFSR_63/R vdd DFFSR_13/D gnd vdd DFFSR
XDFFSR_24 INVX1_16/A DFFSR_9/CLK DFFSR_96/R vdd DFFSR_24/D gnd vdd DFFSR
XDFFSR_46 INVX8_3/A DFFSR_91/CLK DFFSR_9/R vdd DFFSR_46/D gnd vdd DFFSR
XDFFSR_68 DFFSR_68/Q DFFSR_98/CLK DFFSR_93/R vdd DFFSR_68/D gnd vdd DFFSR
XCLKBUF1_33 CLKBUF1_61/Y gnd DFFSR_70/CLK vdd CLKBUF1
XCLKBUF1_22 CLKBUF1_3/A gnd DFFSR_58/CLK vdd CLKBUF1
XDFFSR_57 INVX2_33/A DFFSR_57/CLK DFFSR_63/R vdd DFFSR_57/D gnd vdd DFFSR
XCLKBUF1_11 CLKBUF1_6/A gnd DFFSR_3/CLK vdd CLKBUF1
XDFFSR_79 DFFSR_79/Q DFFSR_4/CLK DFFSR_9/R vdd DFFSR_79/D gnd vdd DFFSR
XCLKBUF1_55 wb_clk_i gnd CLKBUF1_5/A vdd CLKBUF1
XCLKBUF1_44 CLKBUF1_64/Y gnd DFFSR_98/CLK vdd CLKBUF1
XCLKBUF1_66 wb_clk_i gnd CLKBUF1_6/A vdd CLKBUF1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XFILL_20_7_1 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XBUFX4_235 INVX8_11/Y gnd DFFSR_113/S vdd BUFX4
XBUFX4_202 NOR2X1_1/Y gnd BUFX4_202/Y vdd BUFX4
XFILL_18_3_0 gnd vdd FILL
XBUFX4_213 INVX8_8/Y gnd DFFSR_3/R vdd BUFX4
XBUFX4_224 BUFX4_228/A gnd NOR2X1_89/B vdd BUFX4
XBUFX4_257 BUFX4_260/A gnd BUFX4_257/Y vdd BUFX4
XBUFX4_246 BUFX4_250/A gnd BUFX4_246/Y vdd BUFX4
XBUFX4_268 BUFX4_268/A gnd BUFX4_268/Y vdd BUFX4
XNOR2X1_24 NOR3X1_1/B INVX1_79/A gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_35 INVX2_39/A INVX2_40/A gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XNAND3X1_46 OAI21X1_83/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_84/C vdd NAND3X1
XNAND3X1_57 BUFX4_200/Y NAND3X1_57/B AND2X2_3/A gnd NAND3X1_57/Y vdd NAND3X1
XNAND3X1_68 wb_adr_i[2] INVX4_1/Y INVX2_19/Y gnd BUFX4_242/A vdd NAND3X1
XNAND3X1_35 wb_adr_i[4] INVX2_1/Y INVX2_19/Y gnd INVX8_2/A vdd NAND3X1
XNAND3X1_24 AND2X2_3/B OAI21X1_43/Y BUFX4_97/Y gnd OAI21X1_44/C vdd NAND3X1
XNAND3X1_79 NAND3X1_79/A NAND3X1_79/B NAND3X1_79/C gnd DFFSR_88/D vdd NAND3X1
XNAND3X1_13 NAND3X1_9/A OAI21X1_21/Y BUFX4_93/Y gnd OAI21X1_22/C vdd NAND3X1
XNOR2X1_68 INVX4_4/Y XNOR2X1_9/A gnd NOR2X1_70/A vdd NOR2X1
XNOR2X1_57 OR2X2_4/B INVX2_51/Y gnd NOR2X1_60/A vdd NOR2X1
XNOR2X1_79 INVX2_96/A NOR2X1_79/B gnd NOR2X1_79/Y vdd NOR2X1
XNOR2X1_125 INVX2_53/A NOR2X1_99/B gnd OAI22X1_73/B vdd NOR2X1
XNOR2X1_147 INVX2_158/Y NOR2X1_75/B gnd NOR2X1_147/Y vdd NOR2X1
XMUX2X1_20 MUX2X1_38/A MUX2X1_20/B MUX2X1_20/S gnd MUX2X1_20/Y vdd MUX2X1
XNOR2X1_158 BUFX4_125/Y INVX2_156/Y gnd BUFX4_255/A vdd NOR2X1
XMUX2X1_31 wb_dat_i[14] MUX2X1_31/B BUFX4_21/Y gnd MUX2X1_31/Y vdd MUX2X1
XNOR2X1_136 INVX2_110/A BUFX4_176/Y gnd OAI22X1_79/C vdd NOR2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_42/B MUX2X1_42/S gnd MUX2X1_42/Y vdd MUX2X1
XNOR2X1_103 INVX1_31/A NOR2X1_78/B gnd OAI22X1_63/B vdd NOR2X1
XNOR2X1_114 INVX2_62/A NOR2X1_89/B gnd OAI22X1_68/B vdd NOR2X1
XNOR2X1_169 OR2X2_13/B NOR2X1_196/B gnd NOR2X1_169/Y vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XFILL_16_1 gnd vdd FILL
XOAI21X1_609 INVX1_119/Y BUFX4_188/Y OAI21X1_609/C gnd OAI21X1_609/Y vdd OAI21X1
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_7/R vdd DFFSR_1/D gnd vdd DFFSR
XINVX1_27 INVX2_63/A gnd INVX1_27/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XFILL_25_6_1 gnd vdd FILL
XNAND2X1_90 XNOR2X1_4/Y NOR2X1_56/B gnd INVX1_87/A vdd NAND2X1
XFILL_24_1_0 gnd vdd FILL
XFILL_0_6_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_8_7_1 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XNAND3X1_254 INVX4_2/A INVX4_7/A INVX1_124/Y gnd AOI21X1_61/B vdd NAND3X1
XNAND3X1_276 INVX4_4/Y INVX4_3/Y NOR2X1_254/Y gnd NOR2X1_261/A vdd NAND3X1
XNAND3X1_265 INVX4_3/Y AOI21X1_67/A AOI21X1_67/B gnd AOI21X1_68/B vdd NAND3X1
XNAND3X1_210 NOR3X1_4/B OAI21X1_226/Y OAI21X1_227/Y gnd NAND3X1_211/C vdd NAND3X1
XNAND3X1_232 BUFX4_63/Y NAND3X1_232/B NAND3X1_232/C gnd AOI21X1_55/B vdd NAND3X1
XFILL_15_1_0 gnd vdd FILL
XNAND3X1_243 INVX2_147/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_244/C vdd NAND3X1
XNAND3X1_221 INVX2_136/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_223/B vdd NAND3X1
XDFFSR_252 XOR2X1_3/A CLKBUF1_28/Y BUFX4_15/Y vdd DFFSR_252/D gnd vdd DFFSR
XOAI21X1_417 BUFX4_52/Y BUFX4_123/Y NOR2X1_148/Y gnd NOR2X1_191/B vdd OAI21X1
XDFFSR_241 INVX2_86/A CLKBUF1_19/Y BUFX4_8/Y vdd DFFSR_241/D gnd vdd DFFSR
XOAI21X1_406 INVX2_94/Y BUFX4_108/Y OAI21X1_658/C gnd OAI21X1_406/Y vdd OAI21X1
XOAI21X1_428 BUFX4_233/Y OAI21X1_428/B BUFX4_42/Y gnd OAI22X1_86/D vdd OAI21X1
XOAI21X1_439 INVX2_111/Y MUX2X1_29/S OAI21X1_528/C gnd OAI21X1_440/B vdd OAI21X1
XDFFSR_230 INVX2_121/A CLKBUF1_1/Y BUFX4_9/Y vdd DFFSR_230/D gnd vdd DFFSR
XINVX2_81 INVX2_81/A gnd MUX2X1_7/A vdd INVX2
XINVX2_70 INVX2_70/A gnd INVX2_70/Y vdd INVX2
XINVX2_92 INVX2_92/A gnd INVX2_92/Y vdd INVX2
XOAI21X1_11 INVX1_6/Y BUFX4_90/Y NAND2X1_6/Y gnd NAND3X1_8/B vdd OAI21X1
XOAI21X1_66 AND2X2_2/Y INVX2_18/Y OAI21X1_66/C gnd DFFSR_42/D vdd OAI21X1
XOAI21X1_99 INVX2_34/Y BUFX4_20/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_88 AND2X2_2/Y INVX2_28/Y OAI21X1_88/C gnd DFFSR_38/D vdd OAI21X1
XOAI21X1_77 INVX2_23/Y MUX2X1_41/S OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_55 INVX2_13/Y MUX2X1_47/S OAI21X1_83/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_33 INVX2_2/Y BUFX4_20/Y OAI21X1_93/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_44 BUFX4_101/Y INVX2_7/Y OAI21X1_44/C gnd DFFSR_14/D vdd OAI21X1
XOAI21X1_22 BUFX4_102/Y INVX1_11/Y OAI21X1_22/C gnd DFFSR_19/D vdd OAI21X1
XOAI21X1_203 XNOR2X1_5/Y BUFX4_180/Y NAND2X1_91/Y gnd INVX4_5/A vdd OAI21X1
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_236 AOI21X1_63/Y NOR2X1_69/Y OAI21X1_236/C gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_247 INVX2_48/A INVX4_8/Y OAI21X1_247/C gnd OR2X2_9/A vdd OAI21X1
XAND2X2_25 MUX2X1_34/A AND2X2_25/B gnd AND2X2_25/Y vdd AND2X2
XOAI21X1_214 AOI21X1_31/Y AOI21X1_30/Y INVX4_5/Y gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_269 INVX1_35/A NOR2X1_88/B BUFX4_171/Y gnd OAI22X1_55/A vdd OAI21X1
XOAI21X1_258 INVX2_94/A NOR2X1_88/B BUFX4_171/Y gnd OAI22X1_51/A vdd OAI21X1
XOAI21X1_225 AOI21X1_46/Y AOI21X1_47/Y INVX4_5/A gnd OAI21X1_225/Y vdd OAI21X1
XAND2X2_14 AND2X2_14/A BUFX4_266/Y gnd AND2X2_14/Y vdd AND2X2
XNAND2X1_242 BUFX4_6/Y OAI21X1_658/Y gnd OAI21X1_660/C vdd NAND2X1
XNAND2X1_231 BUFX4_2/Y OAI21X1_621/Y gnd OAI21X1_623/C vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_220 INVX4_12/A INVX1_155/Y gnd OAI21X1_570/B vdd NAND2X1
XNAND2X1_253 INVX1_139/A NOR2X1_245/Y gnd OAI21X1_692/B vdd NAND2X1
XFILL_29_0_0 gnd vdd FILL
XFILL_4_0_0 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XDFFSR_36 INVX4_6/A DFFSR_6/CLK DFFSR_80/R vdd DFFSR_36/D gnd vdd DFFSR
XDFFSR_58 INVX2_34/A DFFSR_58/CLK DFFSR_2/R vdd DFFSR_58/D gnd vdd DFFSR
XDFFSR_47 INVX2_39/A DFFSR_2/CLK DFFSR_63/R vdd DFFSR_47/D gnd vdd DFFSR
XDFFSR_14 INVX2_7/A CLKBUF1_8/A DFFSR_7/R vdd DFFSR_14/D gnd vdd DFFSR
XDFFSR_69 DFFSR_69/Q DFFSR_9/CLK DFFSR_96/R vdd DFFSR_69/D gnd vdd DFFSR
XDFFSR_25 INVX1_1/A DFFSR_85/CLK DFFSR_3/R vdd DFFSR_25/D gnd vdd DFFSR
XCLKBUF1_56 wb_clk_i gnd CLKBUF1_2/A vdd CLKBUF1
XCLKBUF1_34 CLKBUF1_5/A gnd DFFSR_55/CLK vdd CLKBUF1
XCLKBUF1_12 CLKBUF1_3/A gnd DFFSR_93/CLK vdd CLKBUF1
XCLKBUF1_23 CLKBUF1_8/A gnd DFFSR_88/CLK vdd CLKBUF1
XCLKBUF1_45 CLKBUF1_63/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_67 wb_clk_i gnd CLKBUF1_3/A vdd CLKBUF1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XINVX1_108 MUX2X1_17/B gnd MUX2X1_18/B vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XBUFX4_236 INVX8_11/Y gnd DFFSR_99/R vdd BUFX4
XBUFX4_269 DFFSR_44/Q gnd BUFX2_80/A vdd BUFX4
XBUFX4_203 BUFX4_207/A gnd NOR2X1_66/B vdd BUFX4
XBUFX4_225 BUFX4_228/A gnd NOR2X1_84/B vdd BUFX4
XBUFX4_247 BUFX4_250/A gnd BUFX4_247/Y vdd BUFX4
XFILL_18_3_1 gnd vdd FILL
XBUFX4_214 INVX8_8/Y gnd DFFSR_96/R vdd BUFX4
XBUFX4_258 BUFX4_260/A gnd BUFX4_258/Y vdd BUFX4
XNAND3X1_14 NAND3X1_9/A OAI21X1_23/Y BUFX4_94/Y gnd OAI21X1_24/C vdd NAND3X1
XNOR2X1_25 OR2X2_2/A OR2X2_2/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_36 INVX2_45/A INVX2_46/A gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_47 INVX2_37/A NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_69 OR2X2_8/B OR2X2_8/A gnd NOR2X1_69/Y vdd NOR2X1
XNAND3X1_36 OAI21X1_65/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_66/C vdd NAND3X1
XNOR2X1_58 INVX2_48/A INVX2_52/Y gnd NOR2X1_62/A vdd NOR2X1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XNAND3X1_47 OAI21X1_85/Y NAND3X1_7/A INVX8_2/Y gnd OAI21X1_86/C vdd NAND3X1
XNAND3X1_69 wb_adr_i[3] INVX4_1/Y INVX2_1/Y gnd BUFX4_135/A vdd NAND3X1
XNAND3X1_25 BUFX4_199/Y OAI21X1_45/Y BUFX4_96/Y gnd OAI21X1_46/C vdd NAND3X1
XNAND3X1_58 BUFX4_199/Y NAND3X1_58/B BUFX4_129/Y gnd NAND3X1_58/Y vdd NAND3X1
XMUX2X1_21 wb_dat_i[28] MUX2X1_21/B BUFX4_92/Y gnd MUX2X1_21/Y vdd MUX2X1
XNOR2X1_126 INVX2_59/A NOR2X1_93/B gnd OAI22X1_74/B vdd NOR2X1
XMUX2X1_10 INVX2_87/Y INVX2_88/Y MUX2X1_8/S gnd MUX2X1_10/Y vdd MUX2X1
XNOR2X1_148 INVX2_159/Y NOR2X1_75/B gnd NOR2X1_148/Y vdd NOR2X1
XNOR2X1_159 INVX2_158/Y INVX2_154/A gnd NOR2X1_159/Y vdd NOR2X1
XMUX2X1_32 MUX2X1_38/A MUX2X1_32/B MUX2X1_32/S gnd MUX2X1_32/Y vdd MUX2X1
XNOR2X1_104 INVX2_137/A BUFX4_176/Y gnd OAI22X1_63/C vdd NOR2X1
XMUX2X1_43 wb_dat_i[0] MUX2X1_43/B MUX2X1_43/S gnd MUX2X1_43/Y vdd MUX2X1
XNOR2X1_137 INVX1_37/A BUFX4_179/Y gnd OAI22X1_79/B vdd NOR2X1
XNOR2X1_115 INVX2_63/A NOR2X1_79/B gnd OAI22X1_68/C vdd NOR2X1
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_2/R vdd DFFSR_2/D gnd vdd DFFSR
XFILL_16_2 gnd vdd FILL
XNAND2X1_80 INVX1_68/Y AND2X2_5/B gnd AND2X2_6/A vdd NAND2X1
XNAND2X1_91 BUFX4_180/Y AND2X2_9/Y gnd NAND2X1_91/Y vdd NAND2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_28 INVX2_65/A gnd INVX1_28/Y vdd INVX1
XINVX1_39 INVX2_78/A gnd INVX1_39/Y vdd INVX1
XFILL_24_1_1 gnd vdd FILL
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XNAND3X1_255 INVX4_6/Y AOI21X1_61/A AOI21X1_61/B gnd AOI21X1_62/B vdd NAND3X1
XNAND3X1_266 INVX2_51/Y INVX1_126/A INVX1_125/Y gnd AOI21X1_69/B vdd NAND3X1
XNAND3X1_222 INVX2_137/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_223/C vdd NAND3X1
XNAND3X1_211 INVX1_86/Y NAND3X1_211/B NAND3X1_211/C gnd NAND3X1_251/B vdd NAND3X1
XNAND3X1_233 INVX2_142/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_235/B vdd NAND3X1
XNAND3X1_200 BUFX4_204/Y NAND3X1_200/B NAND3X1_200/C gnd AOI21X1_50/A vdd NAND3X1
XNAND3X1_244 BUFX4_62/Y NAND3X1_244/B NAND3X1_244/C gnd AOI21X1_57/B vdd NAND3X1
XDFFSR_253 NOR2X1_51/A CLKBUF1_21/Y BUFX4_15/Y vdd DFFSR_253/D gnd vdd DFFSR
XOAI21X1_418 NOR2X1_166/Y MUX2X1_14/B BUFX4_230/Y gnd OAI21X1_418/Y vdd OAI21X1
XOAI21X1_429 BUFX4_52/Y BUFX4_123/Y NOR2X1_151/Y gnd NOR2X1_196/B vdd OAI21X1
XDFFSR_220 INVX1_44/A CLKBUF1_35/Y BUFX4_17/Y vdd DFFSR_220/D gnd vdd DFFSR
XDFFSR_231 INVX2_60/A CLKBUF1_52/Y BUFX4_12/Y vdd DFFSR_231/D gnd vdd DFFSR
XDFFSR_242 INVX2_103/A CLKBUF1_16/Y BUFX4_12/Y vdd DFFSR_242/D gnd vdd DFFSR
XOAI21X1_407 BUFX4_155/Y OAI21X1_407/B OAI21X1_407/C gnd AOI22X1_60/C vdd OAI21X1
XINVX2_82 INVX2_82/A gnd MUX2X1_7/B vdd INVX2
XINVX2_71 INVX2_71/A gnd INVX2_71/Y vdd INVX2
XINVX2_93 INVX2_93/A gnd INVX2_93/Y vdd INVX2
XINVX2_60 INVX2_60/A gnd INVX2_60/Y vdd INVX2
XOAI21X1_34 BUFX4_101/Y INVX2_2/Y OAI21X1_34/C gnd DFFSR_9/D vdd OAI21X1
XOAI21X1_23 INVX1_12/Y NAND2X1_9/B OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_12 OAI21X1_6/A INVX1_6/Y NAND3X1_8/Y gnd DFFSR_30/D vdd OAI21X1
XOAI21X1_45 INVX2_8/Y BUFX4_24/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_67 INVX2_20/Y BUFX4_20/Y OAI21X1_97/C gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_78 AND2X2_2/Y INVX2_23/Y OAI21X1_78/C gnd DFFSR_33/D vdd OAI21X1
XOAI21X1_56 BUFX4_101/Y INVX2_13/Y OAI21X1_56/C gnd DFFSR_4/D vdd OAI21X1
XOAI21X1_89 INVX2_29/Y BUFX4_111/Y OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XOAI21X1_237 OR2X2_7/A OR2X2_7/B INVX4_7/A gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_204 INVX4_7/Y INVX4_6/A XNOR2X1_5/A gnd OAI21X1_205/C vdd OAI21X1
XOAI21X1_215 NOR2X1_64/Y AOI21X1_32/Y OR2X2_6/B gnd BUFX4_61/A vdd OAI21X1
XOAI21X1_226 AOI21X1_48/Y AOI21X1_49/Y INVX4_5/Y gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_248 AND2X2_9/Y INVX4_8/A AOI21X1_74/Y gnd OAI21X1_248/Y vdd OAI21X1
XAND2X2_26 MUX2X1_34/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XOAI21X1_259 INVX2_92/A NOR2X1_89/B BUFX4_80/Y gnd OAI22X1_51/D vdd OAI21X1
XAND2X2_15 AND2X2_15/A BUFX4_268/Y gnd AND2X2_15/Y vdd AND2X2
XFILL_29_0_1 gnd vdd FILL
XNAND2X1_254 BUFX4_4/Y OAI21X1_694/Y gnd OAI21X1_696/C vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_232 INVX8_24/A NOR2X1_226/Y gnd INVX1_156/A vdd NAND2X1
XNAND2X1_210 INVX8_19/A INVX1_146/Y gnd OAI21X1_492/B vdd NAND2X1
XNAND2X1_221 INVX4_12/A AND2X2_20/A gnd OAI21X1_572/B vdd NAND2X1
XNAND2X1_243 INVX8_25/A NOR2X1_226/Y gnd INVX1_157/A vdd NAND2X1
XDFFSR_59 INVX2_35/A CLKBUF1_3/A DFFSR_63/R vdd DFFSR_59/D gnd vdd DFFSR
XDFFSR_37 INVX2_52/A DFFSR_37/CLK DFFSR_80/R vdd DFFSR_37/D gnd vdd DFFSR
XDFFSR_48 INVX2_40/A CLKBUF1_9/Y DFFSR_7/R vdd DFFSR_48/D gnd vdd DFFSR
XDFFSR_26 INVX1_2/A DFFSR_71/CLK DFFSR_7/R vdd DFFSR_26/D gnd vdd DFFSR
XDFFSR_15 INVX2_8/A CLKBUF1_6/A DFFSR_3/R vdd DFFSR_15/D gnd vdd DFFSR
XCLKBUF1_13 CLKBUF1_3/A gnd DFFSR_2/CLK vdd CLKBUF1
XCLKBUF1_46 CLKBUF1_57/Y gnd DFFSR_82/CLK vdd CLKBUF1
XCLKBUF1_57 wb_clk_i gnd CLKBUF1_57/Y vdd CLKBUF1
XCLKBUF1_24 CLKBUF1_6/A gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_35 CLKBUF1_6/A gnd CLKBUF1_35/Y vdd CLKBUF1
XFILL_23_7_0 gnd vdd FILL
XINVX1_109 MUX2X1_31/B gnd MUX2X1_32/B vdd INVX1
XFILL_14_7_0 gnd vdd FILL
XOAI21X1_590 MUX2X1_3/B BUFX4_86/Y OAI21X1_590/C gnd OAI21X1_590/Y vdd OAI21X1
XFILL_4_2 gnd vdd FILL
XBUFX4_237 INVX8_11/Y gnd DFFSR_115/S vdd BUFX4
XBUFX4_226 BUFX4_228/A gnd NOR2X1_88/B vdd BUFX4
XBUFX4_215 INVX8_8/Y gnd DFFSR_2/R vdd BUFX4
XBUFX4_204 BUFX4_207/A gnd BUFX4_204/Y vdd BUFX4
XBUFX4_248 BUFX4_250/A gnd BUFX4_248/Y vdd BUFX4
XBUFX4_259 BUFX4_260/A gnd BUFX4_259/Y vdd BUFX4
XFILL_20_5_0 gnd vdd FILL
XNAND3X1_37 OAI21X1_67/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_68/C vdd NAND3X1
XNAND3X1_48 OAI21X1_87/Y NAND3X1_7/A INVX8_2/Y gnd OAI21X1_88/C vdd NAND3X1
XNAND3X1_15 NAND3X1_9/A OAI21X1_25/Y BUFX4_94/Y gnd OAI21X1_26/C vdd NAND3X1
XNAND3X1_26 BUFX4_199/Y OAI21X1_47/Y BUFX4_96/Y gnd OAI21X1_48/C vdd NAND3X1
XNOR2X1_26 INVX1_70/A NOR2X1_26/B gnd AND2X2_4/A vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNOR2X1_48 OR2X2_5/A OR2X2_5/B gnd NOR2X1_54/A vdd NOR2X1
XNOR2X1_37 INVX2_43/A INVX2_44/A gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_59 NOR3X1_6/A INVX1_89/Y gnd NOR2X1_60/B vdd NOR2X1
XNAND3X1_59 BUFX4_200/Y NAND3X1_59/B BUFX4_130/Y gnd NAND3X1_59/Y vdd NAND3X1
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B gnd NOR2X1_15/Y vdd NOR2X1
XFILL_3_6_0 gnd vdd FILL
XFILL_11_5_0 gnd vdd FILL
XMUX2X1_11 INVX2_89/Y INVX2_90/Y MUX2X1_8/S gnd MUX2X1_11/Y vdd MUX2X1
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_33 wb_dat_i[12] MUX2X1_33/B BUFX4_23/Y gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_22 MUX2X1_34/A MUX2X1_22/B MUX2X1_22/S gnd MUX2X1_22/Y vdd MUX2X1
XNOR2X1_127 INVX2_58/A NOR2X1_93/B gnd OAI22X1_74/C vdd NOR2X1
XNOR2X1_149 NOR2X1_75/A INVX2_155/A gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_116 INVX2_69/A BUFX4_178/Y gnd OAI22X1_69/C vdd NOR2X1
XNOR2X1_105 INVX1_30/A NOR2X1_98/B gnd OAI22X1_64/B vdd NOR2X1
XNOR2X1_138 INVX2_111/A NOR2X1_98/B gnd OAI22X1_80/B vdd NOR2X1
XMUX2X1_44 MUX2X1_48/A MUX2X1_44/B MUX2X1_44/S gnd MUX2X1_44/Y vdd MUX2X1
XFILL_16_3 gnd vdd FILL
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK DFFSR_3/R vdd DFFSR_3/D gnd vdd DFFSR
XINVX1_29 INVX2_64/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_81 AND2X2_4/B XNOR2X1_1/A gnd AND2X2_7/B vdd NAND2X1
XNAND2X1_70 AND2X2_4/A AND2X2_4/B gnd NOR3X1_1/A vdd NAND2X1
XNAND2X1_92 NAND2X1_92/A NAND3X1_91/Y gnd NOR2X1_64/B vdd NAND2X1
XAOI22X1_90 INVX1_158/Y INVX4_10/Y NOR2X1_259/Y AOI22X1_90/D gnd DFFSR_252/D vdd AOI22X1
XNAND3X1_212 INVX2_55/A NAND3X1_212/B NAND3X1_212/C gnd NAND3X1_214/B vdd NAND3X1
XNAND3X1_201 INVX1_114/Y BUFX4_46/Y BUFX4_139/Y gnd NAND3X1_203/B vdd NAND3X1
XNAND3X1_223 BUFX4_204/Y NAND3X1_223/B NAND3X1_223/C gnd AOI21X1_53/A vdd NAND3X1
XNAND3X1_267 AOI21X1_69/B OAI21X1_241/C AND2X2_12/Y gnd OAI21X1_244/A vdd NAND3X1
XNAND3X1_256 INVX4_8/A OAI21X1_235/A OR2X2_5/Y gnd AOI21X1_63/B vdd NAND3X1
XNAND3X1_234 INVX2_143/Y BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_235/C vdd NAND3X1
XNAND3X1_245 INVX2_148/Y BUFX4_74/Y BUFX4_59/Y gnd NAND3X1_247/B vdd NAND3X1
XOAI21X1_419 MUX2X1_14/B BUFX4_92/Y OAI21X1_514/C gnd OAI21X1_420/B vdd OAI21X1
XOAI21X1_408 INVX2_148/Y MUX2X1_37/S OAI21X1_580/C gnd OAI21X1_408/Y vdd OAI21X1
XDFFSR_221 INVX2_83/A CLKBUF1_29/Y BUFX4_8/Y vdd DFFSR_221/D gnd vdd DFFSR
XDFFSR_232 INVX2_136/A CLKBUF1_45/Y BUFX4_12/Y vdd DFFSR_232/D gnd vdd DFFSR
XDFFSR_210 INVX2_105/A CLKBUF1_63/Y BUFX4_12/Y vdd DFFSR_210/D gnd vdd DFFSR
XDFFSR_243 INVX2_68/A CLKBUF1_10/Y BUFX4_12/Y vdd DFFSR_243/D gnd vdd DFFSR
XFILL_25_4_0 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XFILL_8_5_0 gnd vdd FILL
XINVX2_50 XOR2X1_3/A gnd INVX2_50/Y vdd INVX2
XINVX2_83 INVX2_83/A gnd MUX2X1_8/A vdd INVX2
XINVX2_94 INVX2_94/A gnd INVX2_94/Y vdd INVX2
XINVX2_72 INVX2_72/A gnd INVX2_72/Y vdd INVX2
XINVX2_61 INVX2_61/A gnd INVX2_61/Y vdd INVX2
XOAI21X1_68 AND2X2_2/Y INVX2_20/Y OAI21X1_68/C gnd DFFSR_43/D vdd OAI21X1
XFILL_16_4_0 gnd vdd FILL
XOAI21X1_35 INVX2_3/Y BUFX4_22/Y OAI21X1_95/C gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_24 OAI21X1_6/A INVX1_12/Y OAI21X1_24/C gnd DFFSR_20/D vdd OAI21X1
XOAI21X1_13 INVX1_7/Y BUFX4_92/Y NAND2X1_7/Y gnd NAND3X1_9/B vdd OAI21X1
XOAI21X1_57 INVX2_14/Y BUFX4_106/Y OAI21X1_85/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_46 OAI21X1_2/A INVX2_8/Y OAI21X1_46/C gnd DFFSR_15/D vdd OAI21X1
XOAI21X1_79 INVX2_24/Y BUFX4_106/Y OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_238 OR2X2_7/Y INVX4_7/Y INVX2_48/A gnd OAI21X1_238/Y vdd OAI21X1
XOAI21X1_205 INVX4_7/A INVX4_6/Y OAI21X1_205/C gnd XOR2X1_4/A vdd OAI21X1
XOAI21X1_249 INVX4_4/Y XNOR2X1_9/A OAI21X1_249/C gnd AOI21X1_75/B vdd OAI21X1
XOAI21X1_227 AOI21X1_50/Y AOI21X1_51/Y INVX4_5/A gnd OAI21X1_227/Y vdd OAI21X1
XOAI21X1_216 AOI21X1_33/Y AOI21X1_34/Y INVX4_5/A gnd OAI21X1_216/Y vdd OAI21X1
XAND2X2_27 MUX2X1_38/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XNAND2X1_211 INVX8_19/A INVX1_148/Y gnd OAI21X1_504/B vdd NAND2X1
XNAND2X1_200 MUX2X1_41/S wb_dat_i[2] gnd OAI21X1_575/C vdd NAND2X1
XAND2X2_16 AND2X2_16/A BUFX4_268/Y gnd AND2X2_16/Y vdd AND2X2
XNAND2X1_244 NOR2X1_75/Y INVX1_139/A gnd OAI21X1_667/B vdd NAND2X1
XNAND2X1_255 NOR2X1_251/Y MUX2X1_38/A gnd OAI21X1_695/C vdd NAND2X1
XNAND2X1_233 BUFX4_2/Y OAI21X1_624/Y gnd OAI21X1_627/C vdd NAND2X1
XNAND2X1_222 INVX4_12/A NOR2X1_203/Y gnd OAI21X1_574/B vdd NAND2X1
XDFFSR_38 NOR3X1_6/A DFFSR_8/CLK DFFSR_80/R vdd DFFSR_38/D gnd vdd DFFSR
XDFFSR_49 INVX2_41/A DFFSR_4/CLK DFFSR_7/R vdd DFFSR_49/D gnd vdd DFFSR
XDFFSR_27 INVX1_3/A DFFSR_87/CLK DFFSR_96/R vdd DFFSR_27/D gnd vdd DFFSR
XDFFSR_16 INVX2_9/A DFFSR_91/CLK DFFSR_9/R vdd DFFSR_16/D gnd vdd DFFSR
XCLKBUF1_47 CLKBUF1_3/A gnd DFFSR_7/CLK vdd CLKBUF1
XCLKBUF1_25 CLKBUF1_3/A gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_58 wb_clk_i gnd CLKBUF1_8/A vdd CLKBUF1
XCLKBUF1_14 DFFSR_30/CLK gnd DFFSR_92/CLK vdd CLKBUF1
XCLKBUF1_36 DFFSR_30/CLK gnd DFFSR_85/CLK vdd CLKBUF1
XFILL_23_7_1 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XBUFX4_90 wb_sel_i[3] gnd BUFX4_90/Y vdd BUFX4
XFILL_5_3_0 gnd vdd FILL
XFILL_14_7_1 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_591 INVX4_10/A INVX8_22/Y INVX1_152/A gnd NOR2X1_233/B vdd OAI21X1
XOAI21X1_580 INVX2_149/Y BUFX4_108/Y OAI21X1_580/C gnd OAI21X1_580/Y vdd OAI21X1
XFILL_4_3 gnd vdd FILL
XBUFX4_216 INVX8_8/Y gnd DFFSR_63/R vdd BUFX4
XBUFX4_205 BUFX4_207/A gnd BUFX4_205/Y vdd BUFX4
XBUFX4_227 BUFX4_228/A gnd NOR2X1_79/B vdd BUFX4
XBUFX4_238 INVX8_11/Y gnd DFFSR_108/S vdd BUFX4
XBUFX4_249 BUFX4_250/A gnd BUFX4_249/Y vdd BUFX4
XFILL_20_5_1 gnd vdd FILL
XNAND3X1_38 OAI21X1_69/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_70/C vdd NAND3X1
XNAND3X1_49 OAI21X1_89/Y BUFX4_202/Y INVX8_2/Y gnd OAI21X1_90/C vdd NAND3X1
XNAND3X1_27 AND2X2_3/B OAI21X1_49/Y BUFX4_96/Y gnd OAI21X1_50/C vdd NAND3X1
XNAND3X1_16 AND2X2_1/B OAI21X1_27/Y BUFX4_94/Y gnd OAI21X1_28/C vdd NAND3X1
XNOR2X1_27 XNOR2X1_1/B NOR2X1_27/B gnd AND2X2_4/B vdd NOR2X1
XFILL_28_6_1 gnd vdd FILL
XNOR2X1_49 INVX4_7/A NOR2X1_49/B gnd INVX1_88/A vdd NOR2X1
XFILL_27_1_0 gnd vdd FILL
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_16 DFFSR_64/Q NOR2X1_16/B gnd DFFSR_64/D vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XFILL_3_6_1 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B MUX2X1_34/S gnd MUX2X1_34/Y vdd MUX2X1
XFILL_19_6_1 gnd vdd FILL
XMUX2X1_12 MUX2X1_12/A MUX2X1_20/B MUX2X1_8/S gnd MUX2X1_12/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_106 INVX2_138/A NOR2X1_98/B gnd OAI22X1_64/C vdd NOR2X1
XMUX2X1_45 wb_dat_i[31] INVX1_96/A BUFX4_92/Y gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_23 wb_dat_i[26] MUX2X1_23/B BUFX4_87/Y gnd MUX2X1_23/Y vdd MUX2X1
XFILL_16_4 gnd vdd FILL
XNOR2X1_117 INVX2_71/A NOR2X1_87/B gnd OAI22X1_69/B vdd NOR2X1
XNOR2X1_128 INVX2_122/A NOR2X1_96/B gnd OAI22X1_75/C vdd NOR2X1
XNOR2X1_139 INVX1_36/A NOR2X1_71/A gnd OAI22X1_80/C vdd NOR2X1
XDFFSR_4 DFFSR_4/Q DFFSR_4/CLK DFFSR_7/R vdd DFFSR_4/D gnd vdd DFFSR
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_82 INVX1_70/Y AND2X2_5/Y gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_71 NOR2X1_25/Y NOR2X1_29/Y gnd OAI22X1_49/A vdd NAND2X1
XNAND2X1_60 MUX2X1_25/B BUFX4_117/Y gnd NAND3X1_81/A vdd NAND2X1
XNAND2X1_93 XOR2X1_4/B XOR2X1_4/A gnd NAND2X1_93/Y vdd NAND2X1
XAOI21X1_220 INVX2_76/Y OAI21X1_692/B BUFX4_265/Y gnd OAI21X1_692/C vdd AOI21X1
XAOI22X1_80 INVX2_125/Y BUFX4_3/Y AOI22X1_80/C AOI22X1_80/D gnd DFFSR_150/D vdd AOI22X1
XNAND3X1_257 INVX4_3/A AOI21X1_63/A AOI21X1_63/B gnd OAI21X1_236/C vdd NAND3X1
XNAND3X1_213 NAND3X1_213/A NAND3X1_213/B INVX2_55/Y gnd NAND3X1_214/C vdd NAND3X1
XNAND3X1_235 BUFX4_207/Y NAND3X1_235/B NAND3X1_235/C gnd AOI21X1_56/A vdd NAND3X1
XNAND3X1_224 INVX1_119/Y BUFX4_51/Y BUFX4_140/Y gnd NAND3X1_226/B vdd NAND3X1
XNAND3X1_202 INVX2_123/Y BUFX4_73/Y BUFX4_56/Y gnd NAND3X1_203/C vdd NAND3X1
XNAND3X1_246 INVX2_149/Y BUFX4_47/Y BUFX4_136/Y gnd NAND3X1_247/C vdd NAND3X1
XNAND3X1_268 AOI21X1_62/B AND2X2_12/Y OAI21X1_243/Y gnd NAND3X1_272/C vdd NAND3X1
XFILL_14_1 gnd vdd FILL
XDFFSR_200 INVX2_138/A CLKBUF1_1/Y BUFX4_9/Y vdd DFFSR_200/D gnd vdd DFFSR
XOAI21X1_409 BUFX4_54/Y BUFX4_126/Y INVX1_140/A gnd INVX1_145/A vdd OAI21X1
XDFFSR_244 BUFX2_1/A CLKBUF1_5/Y BUFX4_14/Y vdd DFFSR_244/D gnd vdd DFFSR
XDFFSR_222 INVX1_50/A CLKBUF1_25/Y BUFX4_16/Y vdd DFFSR_222/D gnd vdd DFFSR
XDFFSR_233 INVX2_97/A CLKBUF1_41/Y BUFX4_9/Y vdd DFFSR_233/D gnd vdd DFFSR
XDFFSR_211 INVX2_67/A CLKBUF1_19/Y BUFX4_10/Y vdd DFFSR_211/D gnd vdd DFFSR
XFILL_25_4_1 gnd vdd FILL
XFILL_0_4_1 gnd vdd FILL
XINVX2_51 NOR3X1_6/A gnd INVX2_51/Y vdd INVX2
XINVX2_40 INVX2_40/A gnd INVX2_40/Y vdd INVX2
XINVX2_73 INVX2_73/A gnd INVX2_73/Y vdd INVX2
XFILL_7_0_0 gnd vdd FILL
XFILL_8_5_1 gnd vdd FILL
XINVX2_62 INVX2_62/A gnd INVX2_62/Y vdd INVX2
XINVX2_84 INVX2_84/A gnd MUX2X1_8/B vdd INVX2
XFILL_16_4_1 gnd vdd FILL
XINVX2_95 INVX2_95/A gnd INVX2_95/Y vdd INVX2
XOAI21X1_69 INVX2_21/Y BUFX4_21/Y OAI21X1_99/C gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_25 INVX1_13/Y MUX2X1_29/S OAI21X1_25/C gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_14 OAI21X1_6/A INVX1_7/Y NAND3X1_9/Y gnd DFFSR_31/D vdd OAI21X1
XOAI21X1_58 OAI21X1_2/A INVX2_14/Y OAI21X1_58/C gnd DFFSR_5/D vdd OAI21X1
XOAI21X1_36 OAI21X1_2/A INVX2_3/Y OAI21X1_36/C gnd DFFSR_10/D vdd OAI21X1
XOAI21X1_47 INVX2_9/Y BUFX4_26/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_239 OR2X2_7/Y INVX4_7/Y INVX2_48/Y gnd OAI21X1_239/Y vdd OAI21X1
XOAI21X1_217 AOI21X1_35/Y AOI21X1_36/Y INVX8_13/Y gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_228 AOI21X1_52/Y AOI21X1_53/Y INVX4_5/A gnd AOI21X1_54/B vdd OAI21X1
XOAI21X1_206 NOR2X1_63/Y AOI21X1_29/Y OR2X2_6/B gnd BUFX4_142/A vdd OAI21X1
XAND2X2_28 MUX2X1_34/A AND2X2_28/B gnd AND2X2_28/Y vdd AND2X2
XNAND2X1_201 NOR2X1_159/Y INVX1_139/A gnd OAI21X1_405/B vdd NAND2X1
XNAND2X1_212 INVX4_11/A NOR2X1_195/Y gnd OAI21X1_519/B vdd NAND2X1
XNAND2X1_234 NOR2X1_228/Y MUX2X1_42/A gnd OAI21X1_626/C vdd NAND2X1
XAND2X2_17 AND2X2_17/A INVX4_11/A gnd AND2X2_17/Y vdd AND2X2
XNAND2X1_223 INVX4_12/A NOR2X1_205/Y gnd OAI21X1_579/B vdd NAND2X1
XNAND2X1_245 BUFX4_20/Y wb_dat_i[15] gnd OAI21X1_694/C vdd NAND2X1
XNAND2X1_256 BUFX4_1/Y OAI21X1_697/Y gnd OAI21X1_700/C vdd NAND2X1
XDFFSR_28 INVX1_4/A DFFSR_88/CLK DFFSR_7/R vdd DFFSR_28/D gnd vdd DFFSR
XDFFSR_17 INVX1_9/A DFFSR_92/CLK DFFSR_95/R vdd DFFSR_17/D gnd vdd DFFSR
XDFFSR_39 XOR2X1_3/B DFFSR_99/CLK DFFSR_93/R vdd DFFSR_39/D gnd vdd DFFSR
XCLKBUF1_15 CLKBUF1_6/A gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_37 CLKBUF1_2/A gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_48 CLKBUF1_2/A gnd DFFSR_37/CLK vdd CLKBUF1
XCLKBUF1_26 CLKBUF1_64/Y gnd DFFSR_57/CLK vdd CLKBUF1
XBUFX4_91 wb_sel_i[3] gnd BUFX4_91/Y vdd BUFX4
XCLKBUF1_59 wb_clk_i gnd CLKBUF1_4/A vdd CLKBUF1
XBUFX4_80 NOR3X1_8/Y gnd BUFX4_80/Y vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 XNOR2X1_1/A XNOR2X1_1/B gnd XNOR2X1_1/Y vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XOAI21X1_592 AND2X2_21/B INVX1_93/A BUFX4_162/Y gnd OAI21X1_593/B vdd OAI21X1
XOAI21X1_581 BUFX4_127/Y INVX8_22/Y AND2X2_17/A gnd NOR2X1_230/B vdd OAI21X1
XOAI21X1_570 BUFX4_159/Y OAI21X1_570/B OAI21X1_570/C gnd AOI22X1_78/C vdd OAI21X1
XFILL_4_4 gnd vdd FILL
XBUFX4_228 BUFX4_228/A gnd NOR2X1_93/B vdd BUFX4
XBUFX4_217 BUFX4_220/A gnd INVX8_4/A vdd BUFX4
XBUFX4_239 BUFX4_242/A gnd OAI22X1_7/A vdd BUFX4
XBUFX4_206 BUFX4_207/A gnd BUFX4_206/Y vdd BUFX4
XAND2X2_1 BUFX4_95/Y AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_28 NOR2X1_28/A INVX1_68/A gnd AND2X2_5/A vdd NOR2X1
XNAND3X1_39 OAI21X1_71/Y AND2X2_2/B INVX8_2/Y gnd OAI21X1_72/C vdd NAND3X1
XNAND3X1_28 BUFX4_200/Y OAI21X1_51/Y BUFX4_97/Y gnd OAI21X1_52/C vdd NAND3X1
XNOR2X1_17 NOR2X1_1/B NOR2X1_17/B gnd INVX8_20/A vdd NOR2X1
XNAND3X1_17 NAND3X1_9/A OAI21X1_29/Y BUFX4_94/Y gnd OAI21X1_30/C vdd NAND3X1
XNOR2X1_39 XOR2X1_1/A XOR2X1_1/B gnd AND2X2_5/B vdd NOR2X1
XFILL_27_1_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_13 MUX2X1_13/A MUX2X1_13/B MUX2X1_9/S gnd MUX2X1_13/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XNOR2X1_107 INVX1_43/A NOR2X1_82/B gnd OAI22X1_65/B vdd NOR2X1
XNOR2X1_118 INVX2_67/A NOR2X1_79/B gnd OAI22X1_70/B vdd NOR2X1
XNOR2X1_129 INVX1_25/A NOR2X1_96/B gnd OAI22X1_75/B vdd NOR2X1
XMUX2X1_35 wb_dat_i[6] MUX2X1_35/B MUX2X1_35/S gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_46 MUX2X1_48/A INVX1_96/Y MUX2X1_46/S gnd MUX2X1_46/Y vdd MUX2X1
XMUX2X1_24 MUX2X1_48/A MUX2X1_24/B MUX2X1_24/S gnd MUX2X1_24/Y vdd MUX2X1
XDFFSR_5 DFFSR_5/Q DFFSR_5/CLK DFFSR_9/R vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_50 NAND2X1_50/A NAND2X1_50/B gnd DFFSR_80/D vdd NAND2X1
XNAND2X1_61 MUX2X1_23/B BUFX4_114/Y gnd NAND3X1_82/A vdd NAND2X1
XNAND2X1_94 NAND2X1_94/A OR2X2_4/Y gnd INVX1_91/A vdd NAND2X1
XNAND2X1_72 INVX1_66/Y INVX1_67/Y gnd NOR2X1_33/A vdd NAND2X1
XNAND2X1_83 NAND2X1_83/A NAND2X1_83/B gnd DFFSR_111/D vdd NAND2X1
XAOI21X1_210 BUFX4_259/Y OAI21X1_672/Y BUFX4_5/Y gnd AOI22X1_84/D vdd AOI21X1
XAOI21X1_221 BUFX4_265/Y OAI21X1_693/Y BUFX4_246/Y gnd AOI22X1_89/D vdd AOI21X1
XAOI22X1_81 INVX2_149/Y BUFX4_3/Y AOI22X1_81/C AOI22X1_81/D gnd DFFSR_148/D vdd AOI22X1
XAOI22X1_70 INVX2_116/Y BUFX4_5/Y AOI22X1_70/C AOI22X1_70/D gnd DFFSR_174/D vdd AOI22X1
XNAND3X1_269 INVX1_129/A INVX2_151/A NAND3X1_272/C gnd AOI21X1_73/A vdd NAND3X1
XNAND3X1_258 INVX4_6/A AOI21X1_61/A AOI21X1_61/B gnd NAND3X1_258/Y vdd NAND3X1
XNAND3X1_214 INVX4_5/Y NAND3X1_214/B NAND3X1_214/C gnd AOI21X1_54/A vdd NAND3X1
XNAND3X1_236 INVX1_121/Y BUFX4_49/Y BUFX4_142/Y gnd NAND3X1_238/B vdd NAND3X1
XNAND3X1_203 BUFX4_62/Y NAND3X1_203/B NAND3X1_203/C gnd AOI21X1_50/B vdd NAND3X1
XNAND3X1_225 INVX2_138/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_226/C vdd NAND3X1
XNAND3X1_247 BUFX4_205/Y NAND3X1_247/B NAND3X1_247/C gnd AOI21X1_58/A vdd NAND3X1
XDFFSR_223 INVX2_56/A CLKBUF1_21/Y BUFX4_8/Y vdd DFFSR_223/D gnd vdd DFFSR
XFILL_14_2 gnd vdd FILL
XDFFSR_201 INVX2_99/A CLKBUF1_52/Y BUFX4_16/Y vdd DFFSR_201/D gnd vdd DFFSR
XDFFSR_212 INVX1_20/A CLKBUF1_16/Y BUFX4_9/Y vdd DFFSR_212/D gnd vdd DFFSR
XDFFSR_234 INVX2_109/A CLKBUF1_40/Y BUFX4_16/Y vdd DFFSR_234/D gnd vdd DFFSR
XDFFSR_245 DFFSR_245/Q CLKBUF1_2/Y BUFX4_14/Y vdd DFFSR_245/D gnd vdd DFFSR
XINVX2_52 INVX2_52/A gnd INVX2_52/Y vdd INVX2
XINVX2_85 INVX2_85/A gnd MUX2X1_9/A vdd INVX2
XINVX2_30 INVX2_30/A gnd INVX2_30/Y vdd INVX2
XINVX2_96 INVX2_96/A gnd INVX2_96/Y vdd INVX2
XINVX2_74 INVX2_74/A gnd INVX2_74/Y vdd INVX2
XFILL_7_0_1 gnd vdd FILL
XINVX2_41 INVX2_41/A gnd INVX2_41/Y vdd INVX2
XINVX2_63 INVX2_63/A gnd INVX2_63/Y vdd INVX2
XOAI21X1_37 INVX2_4/Y BUFX4_24/Y OAI21X1_97/C gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_59 INVX2_15/Y BUFX4_108/Y OAI21X1_87/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_26 BUFX4_102/Y INVX1_13/Y OAI21X1_26/C gnd DFFSR_21/D vdd OAI21X1
XOAI21X1_15 INVX1_8/Y BUFX4_87/Y NAND2X1_8/Y gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_48 OAI21X1_2/A INVX2_9/Y OAI21X1_48/C gnd DFFSR_16/D vdd OAI21X1
XOAI21X1_207 OR2X2_6/B OR2X2_6/A BUFX4_142/Y gnd INVX2_55/A vdd OAI21X1
XAND2X2_29 MUX2X1_38/A AND2X2_29/B gnd AND2X2_29/Y vdd AND2X2
XOAI21X1_229 AOI21X1_55/Y AOI21X1_56/Y INVX4_5/Y gnd AOI21X1_59/A vdd OAI21X1
XOAI21X1_218 AOI21X1_37/Y AOI21X1_38/Y INVX8_13/A gnd OAI21X1_218/Y vdd OAI21X1
XAND2X2_18 AND2X2_18/A INVX4_11/A gnd AND2X2_18/Y vdd AND2X2
XNAND2X1_224 BUFX4_6/Y OAI21X1_590/Y gnd OAI21X1_593/C vdd NAND2X1
XNAND2X1_235 BUFX4_6/Y OAI21X1_630/Y gnd OAI21X1_632/C vdd NAND2X1
XNAND2X1_202 MUX2X1_43/S wb_dat_i[1] gnd OAI21X1_658/C vdd NAND2X1
XNAND2X1_257 NOR2X1_252/Y INVX8_14/A gnd OAI21X1_699/C vdd NAND2X1
XNAND2X1_213 INVX4_11/A INVX1_155/Y gnd OAI21X1_534/B vdd NAND2X1
XNAND2X1_246 NOR2X1_71/Y NOR2X1_245/Y gnd OAI21X1_669/B vdd NAND2X1
XFILL_26_7_0 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XFILL_17_7_0 gnd vdd FILL
XDFFSR_29 INVX1_5/A CLKBUF1_3/A DFFSR_80/R vdd DFFSR_29/D gnd vdd DFFSR
XDFFSR_18 INVX1_10/A DFFSR_3/CLK DFFSR_95/R vdd DFFSR_18/D gnd vdd DFFSR
XCLKBUF1_27 CLKBUF1_57/Y gnd DFFSR_87/CLK vdd CLKBUF1
XCLKBUF1_38 CLKBUF1_4/A gnd DFFSR_9/CLK vdd CLKBUF1
XCLKBUF1_16 CLKBUF1_54/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_49 CLKBUF1_2/A gnd CLKBUF1_49/Y vdd CLKBUF1
XBUFX4_92 wb_sel_i[3] gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 BUFX4_85/A gnd BUFX4_81/Y vdd BUFX4
XBUFX4_70 INVX8_5/Y gnd BUFX4_70/Y vdd BUFX4
XXNOR2X1_2 NOR3X1_3/C INVX2_47/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XOAI21X1_560 NOR2X1_210/Y MUX2X1_6/A BUFX4_148/Y gnd OAI21X1_560/Y vdd OAI21X1
XOAI21X1_593 AND2X2_21/Y OAI21X1_593/B OAI21X1_593/C gnd DFFSR_143/D vdd OAI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_582 BUFX4_124/Y INVX8_20/Y MUX2X1_18/Y gnd OAI21X1_583/C vdd OAI21X1
XOAI21X1_571 INVX2_134/Y MUX2X1_47/S OAI21X1_651/C gnd OAI21X1_571/Y vdd OAI21X1
XFILL_23_5_0 gnd vdd FILL
XBUFX4_207 BUFX4_207/A gnd BUFX4_207/Y vdd BUFX4
XBUFX4_218 BUFX4_220/A gnd OAI22X1_5/D vdd BUFX4
XBUFX4_229 INVX8_18/Y gnd BUFX4_229/Y vdd BUFX4
XFILL_6_6_0 gnd vdd FILL
XFILL_14_5_0 gnd vdd FILL
XAND2X2_2 INVX8_2/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XOAI21X1_390 OAI21X1_390/A BUFX4_245/Y OAI21X1_390/C gnd DFFSR_222/D vdd OAI21X1
XFILL_2_2 gnd vdd FILL
XNOR2X1_29 NOR3X1_1/A NOR2X1_29/B gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_18 NOR2X1_1/B NOR2X1_18/B gnd INVX8_22/A vdd NOR2X1
XNAND3X1_18 NAND3X1_9/A OAI21X1_31/Y BUFX4_94/Y gnd OAI21X1_32/C vdd NAND3X1
XNAND3X1_29 AND2X2_1/B OAI21X1_53/Y BUFX4_95/Y gnd OAI21X1_54/C vdd NAND3X1
XMUX2X1_25 wb_dat_i[25] MUX2X1_25/B BUFX4_88/Y gnd MUX2X1_26/B vdd MUX2X1
XMUX2X1_14 MUX2X1_14/A MUX2X1_14/B MUX2X1_9/S gnd MUX2X1_14/Y vdd MUX2X1
XNOR2X1_108 INVX2_140/A NOR2X1_82/B gnd OAI22X1_65/C vdd NOR2X1
XNOR2X1_119 INVX2_70/A NOR2X1_79/B gnd OAI22X1_70/C vdd NOR2X1
XMUX2X1_47 wb_dat_i[7] INVX1_99/A MUX2X1_47/S gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_36 MUX2X1_48/A MUX2X1_36/B MUX2X1_36/S gnd MUX2X1_36/Y vdd MUX2X1
XDFFSR_6 DFFSR_6/Q DFFSR_6/CLK DFFSR_7/R vdd DFFSR_6/D gnd vdd DFFSR
XNAND2X1_84 INVX1_75/A NOR3X1_1/Y gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_73 NOR2X1_34/Y NOR2X1_35/Y gnd NOR2X1_38/A vdd NAND2X1
XNAND2X1_95 BUFX4_180/Y INVX1_91/A gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_62 INVX1_93/A BUFX4_117/Y gnd NAND3X1_83/A vdd NAND2X1
XNAND2X1_40 AOI21X1_6/Y NOR2X1_7/Y gnd DFFSR_70/D vdd NAND2X1
XNAND2X1_51 INVX1_122/A BUFX4_116/Y gnd NAND3X1_72/A vdd NAND2X1
XAOI21X1_200 BUFX4_260/Y OAI21X1_575/Y BUFX4_3/Y gnd AOI22X1_80/D vdd AOI21X1
XAOI21X1_222 BUFX4_123/Y XNOR2X1_14/Y NOR2X1_254/Y gnd DFFSR_246/D vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XAOI21X1_211 NOR2X1_247/Y BUFX4_160/Y OAI21X1_673/Y gnd OAI22X1_119/C vdd AOI21X1
XAOI22X1_82 INVX2_72/Y BUFX4_247/Y AOI22X1_82/C AOI22X1_82/D gnd DFFSR_227/D vdd AOI22X1
XAOI22X1_71 INVX2_137/Y BUFX4_1/Y AOI22X1_71/C AOI22X1_71/D gnd DFFSR_168/D vdd AOI22X1
XAOI22X1_60 INVX2_148/Y BUFX4_245/Y AOI22X1_60/C AOI22X1_60/D gnd DFFSR_212/D vdd
+ AOI22X1
XFILL_28_4_0 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XNAND3X1_259 INVX4_2/A INVX4_7/Y INVX1_124/Y gnd NAND3X1_260/C vdd NAND3X1
XNAND3X1_237 INVX2_144/Y BUFX4_75/Y BUFX4_58/Y gnd NAND3X1_238/C vdd NAND3X1
XNAND3X1_226 BUFX4_62/Y NAND3X1_226/B NAND3X1_226/C gnd AOI21X1_53/B vdd NAND3X1
XNAND3X1_215 INVX2_133/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_217/B vdd NAND3X1
XNAND3X1_204 INVX2_124/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_206/B vdd NAND3X1
XNAND3X1_248 MUX2X1_44/B BUFX4_47/Y BUFX4_136/Y gnd NAND3X1_250/B vdd NAND3X1
XFILL_11_3_0 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XDFFSR_246 OR2X2_5/A CLKBUF1_49/Y BUFX4_15/Y vdd DFFSR_246/D gnd vdd DFFSR
XDFFSR_224 INVX1_56/A CLKBUF1_60/Y BUFX4_8/Y vdd DFFSR_224/D gnd vdd DFFSR
XDFFSR_213 INVX2_94/A CLKBUF1_9/Y BUFX4_10/Y vdd DFFSR_213/D gnd vdd DFFSR
XDFFSR_202 INVX2_111/A CLKBUF1_45/Y BUFX4_12/Y vdd DFFSR_202/D gnd vdd DFFSR
XDFFSR_235 INVX2_73/A CLKBUF1_35/Y BUFX4_16/Y vdd DFFSR_235/D gnd vdd DFFSR
XINVX2_53 INVX2_53/A gnd MUX2X1_2/A vdd INVX2
XINVX2_20 MUX2X1_1/S gnd INVX2_20/Y vdd INVX2
XINVX2_42 INVX2_42/A gnd INVX2_42/Y vdd INVX2
XINVX2_31 INVX2_31/A gnd INVX2_31/Y vdd INVX2
XINVX2_86 INVX2_86/A gnd MUX2X1_9/B vdd INVX2
XINVX2_75 INVX2_75/A gnd INVX2_75/Y vdd INVX2
XINVX2_97 INVX2_97/A gnd INVX2_97/Y vdd INVX2
XINVX2_64 INVX2_64/A gnd INVX2_64/Y vdd INVX2
XOAI21X1_16 OAI21X1_6/A INVX1_8/Y OAI21X1_16/C gnd DFFSR_32/D vdd OAI21X1
XOAI21X1_38 BUFX4_101/Y INVX2_4/Y OAI21X1_38/C gnd DFFSR_11/D vdd OAI21X1
XOAI21X1_49 INVX2_10/Y BUFX4_106/Y OAI21X1_77/C gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_27 INVX1_14/Y BUFX4_188/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_208 INVX2_48/A INVX2_52/Y NAND2X1_93/Y gnd XOR2X1_5/A vdd OAI21X1
XOAI21X1_219 AOI21X1_39/Y AOI21X1_40/Y INVX4_5/A gnd OAI21X1_219/Y vdd OAI21X1
XAND2X2_19 AND2X2_19/A INVX4_11/A gnd AND2X2_19/Y vdd AND2X2
XNAND2X1_258 INVX4_9/A AND2X2_9/Y gnd OAI21X1_705/C vdd NAND2X1
XNAND2X1_225 NOR2X1_219/Y MUX2X1_34/A gnd OAI21X1_598/C vdd NAND2X1
XNAND2X1_236 BUFX4_6/Y OAI21X1_635/Y gnd OAI21X1_637/C vdd NAND2X1
XNAND2X1_214 INVX4_11/A NOR2X1_203/Y gnd OAI21X1_539/B vdd NAND2X1
XNAND2X1_247 MUX2X1_29/S wb_dat_i[23] gnd OAI21X1_697/C vdd NAND2X1
XNAND2X1_203 NOR2X1_160/Y INVX1_139/A gnd OAI21X1_407/B vdd NAND2X1
XFILL_26_7_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XFILL_17_7_1 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XDFFSR_19 INVX1_11/A CLKBUF1_6/Y DFFSR_95/R vdd DFFSR_19/D gnd vdd DFFSR
XCLKBUF1_28 CLKBUF1_61/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_39 CLKBUF1_3/A gnd DFFSR_99/CLK vdd CLKBUF1
XCLKBUF1_17 CLKBUF1_57/Y gnd DFFSR_91/CLK vdd CLKBUF1
XBUFX4_82 BUFX4_85/A gnd MUX2X1_8/S vdd BUFX4
XBUFX4_93 INVX8_1/Y gnd BUFX4_93/Y vdd BUFX4
XBUFX4_71 BUFX4_76/A gnd BUFX4_71/Y vdd BUFX4
XBUFX4_60 BUFX4_61/A gnd BUFX4_60/Y vdd BUFX4
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_3/A vdd OR2X2
XXNOR2X1_3 OR2X2_5/B INVX4_3/A gnd XNOR2X1_3/Y vdd XNOR2X1
XOAI21X1_561 MUX2X1_6/A BUFX4_19/Y OAI21X1_641/C gnd OAI21X1_562/B vdd OAI21X1
XOAI21X1_550 INVX2_89/Y BUFX4_23/Y OAI21X1_630/C gnd OAI21X1_551/B vdd OAI21X1
XOAI21X1_594 BUFX4_121/Y INVX8_22/Y NOR2X1_195/Y gnd NOR2X1_234/B vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_583 BUFX4_161/Y MUX2X1_17/Y OAI21X1_583/C gnd DFFSR_146/D vdd OAI21X1
XOAI21X1_572 BUFX4_159/Y OAI21X1_572/B OAI21X1_572/C gnd AOI22X1_79/C vdd OAI21X1
XFILL_23_5_1 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XBUFX4_219 BUFX4_220/A gnd OAI22X1_8/D vdd BUFX4
XBUFX4_208 INVX8_8/Y gnd DFFSR_7/R vdd BUFX4
XFILL_5_1_0 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XOAI21X1_391 BUFX4_156/Y OAI21X1_391/B OAI21X1_391/C gnd AOI22X1_52/C vdd OAI21X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_380 BUFX4_144/Y BUFX4_255/Y INVX2_106/A gnd OAI21X1_381/C vdd OAI21X1
XNAND3X1_19 BUFX4_199/Y OAI21X1_33/Y BUFX4_96/Y gnd OAI21X1_34/C vdd NAND3X1
XNOR2X1_19 NOR2X1_1/B INVX8_7/A gnd NOR2X1_19/Y vdd NOR2X1
XMUX2X1_26 MUX2X1_26/A MUX2X1_26/B MUX2X1_26/S gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_15 MUX2X1_15/A MUX2X1_15/B MUX2X1_6/S gnd MUX2X1_15/Y vdd MUX2X1
XNOR2X1_109 INVX1_42/A NOR2X1_88/B gnd OAI22X1_66/B vdd NOR2X1
XMUX2X1_37 wb_dat_i[5] MUX2X1_37/B MUX2X1_37/S gnd MUX2X1_37/Y vdd MUX2X1
XMUX2X1_48 MUX2X1_48/A INVX1_99/Y MUX2X1_48/S gnd MUX2X1_48/Y vdd MUX2X1
XDFFSR_7 DFFSR_7/Q DFFSR_7/CLK DFFSR_7/R vdd DFFSR_7/D gnd vdd DFFSR
XNAND2X1_74 NOR2X1_36/Y NOR2X1_37/Y gnd NOR2X1_38/B vdd NAND2X1
XNAND2X1_85 NAND2X1_85/A NAND2X1_85/B gnd DFFSR_113/D vdd NAND2X1
XNAND2X1_96 BUFX4_180/Y AND2X2_10/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_63 MUX2X1_21/B BUFX4_117/Y gnd NAND3X1_84/A vdd NAND2X1
XNAND2X1_30 MUX2X1_43/S wb_dat_i[5] gnd OAI21X1_87/C vdd NAND2X1
XNAND2X1_52 INVX1_103/A BUFX4_116/Y gnd NAND3X1_73/A vdd NAND2X1
XNAND2X1_41 AOI21X1_7/Y NOR2X1_8/Y gnd DFFSR_71/D vdd NAND2X1
XAOI21X1_223 NOR2X1_262/Y NOR2X1_259/B NOR2X1_261/Y gnd OAI21X1_711/C vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_201 NOR2X1_212/Y BUFX4_154/Y OAI21X1_576/Y gnd OAI22X1_117/C vdd AOI21X1
XAOI21X1_212 INVX2_75/Y OR2X2_13/Y BUFX4_251/Y gnd OAI21X1_677/C vdd AOI21X1
XAOI22X1_50 MUX2X1_13/A BUFX4_250/Y AOI22X1_50/C AOI22X1_50/D gnd DFFSR_224/D vdd
+ AOI22X1
XAOI22X1_72 INVX2_122/Y BUFX4_1/Y AOI22X1_72/C AOI22X1_72/D gnd DFFSR_166/D vdd AOI22X1
XAOI22X1_61 INVX2_105/Y BUFX4_145/Y AOI22X1_61/C AOI22X1_61/D gnd DFFSR_210/D vdd
+ AOI22X1
XAOI22X1_83 INVX2_73/Y BUFX4_248/Y AOI22X1_83/C AOI22X1_83/D gnd DFFSR_235/D vdd AOI22X1
XFILL_28_4_1 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XNAND3X1_205 INVX2_125/Y BUFX4_47/Y BUFX4_141/Y gnd NAND3X1_206/C vdd NAND3X1
XNAND3X1_238 BUFX4_63/Y NAND3X1_238/B NAND3X1_238/C gnd AOI21X1_56/B vdd NAND3X1
XNAND3X1_227 INVX2_139/Y BUFX4_76/Y BUFX4_57/Y gnd NAND3X1_229/B vdd NAND3X1
XNAND3X1_216 INVX2_134/Y BUFX4_47/Y BUFX4_139/Y gnd NAND3X1_217/C vdd NAND3X1
XNAND3X1_249 INVX2_150/Y BUFX4_72/Y BUFX4_60/Y gnd NAND3X1_250/C vdd NAND3X1
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 OAI22X1_7/A INVX1_19/Y INVX1_18/Y OAI22X1_7/D gnd NOR2X1_2/B vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XDFFSR_247 OR2X2_5/B DFFSR_37/CLK BUFX4_15/Y vdd DFFSR_247/D gnd vdd DFFSR
XDFFSR_225 INVX2_85/A CLKBUF1_54/Y BUFX4_17/Y vdd DFFSR_225/D gnd vdd DFFSR
XDFFSR_203 INVX2_75/A DFFSR_83/CLK BUFX4_13/Y vdd DFFSR_203/D gnd vdd DFFSR
XDFFSR_214 INVX1_26/A CLKBUF1_7/Y BUFX4_9/Y vdd DFFSR_214/D gnd vdd DFFSR
XDFFSR_236 INVX2_139/A DFFSR_86/CLK BUFX4_10/Y vdd DFFSR_236/D gnd vdd DFFSR
XINVX2_21 OR2X2_9/B gnd INVX2_21/Y vdd INVX2
XINVX2_10 DFFSR_1/Q gnd INVX2_10/Y vdd INVX2
XINVX2_54 INVX2_54/A gnd MUX2X1_2/B vdd INVX2
XINVX2_87 INVX2_87/A gnd INVX2_87/Y vdd INVX2
XINVX2_32 INVX2_32/A gnd INVX2_32/Y vdd INVX2
XINVX2_98 INVX2_98/A gnd INVX2_98/Y vdd INVX2
XINVX2_65 INVX2_65/A gnd INVX2_65/Y vdd INVX2
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XINVX2_76 INVX2_76/A gnd INVX2_76/Y vdd INVX2
XOAI21X1_28 OAI21X1_6/A INVX1_14/Y OAI21X1_28/C gnd DFFSR_22/D vdd OAI21X1
XOAI21X1_17 INVX1_9/Y BUFX4_185/Y NAND2X1_9/Y gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_39 INVX2_5/Y BUFX4_26/Y OAI21X1_99/C gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_209 INVX1_88/Y INVX2_48/A OR2X2_4/B gnd NAND2X1_94/A vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XNAND2X1_259 INVX4_6/A INVX4_10/Y gnd OAI21X1_706/C vdd NAND2X1
XNAND2X1_237 BUFX4_6/Y OAI21X1_638/Y gnd OAI21X1_640/C vdd NAND2X1
XNAND2X1_248 INVX4_11/A NOR2X1_246/Y gnd OAI21X1_671/B vdd NAND2X1
XNAND2X1_226 BUFX4_2/Y OAI21X1_605/Y gnd OAI21X1_608/C vdd NAND2X1
XNAND2X1_215 INVX4_11/A NOR2X1_205/Y gnd OAI21X1_545/B vdd NAND2X1
XNAND2X1_204 MUX2X1_35/S wb_dat_i[0] gnd OAI21X1_580/C vdd NAND2X1
XFILL_25_2_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XOAI21X1_710 OR2X2_4/Y INVX4_9/Y XOR2X1_3/A gnd AOI22X1_90/D vdd OAI21X1
XFILL_8_3_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XCLKBUF1_29 CLKBUF1_61/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XCLKBUF1_18 CLKBUF1_64/Y gnd DFFSR_1/CLK vdd CLKBUF1
XBUFX4_50 OR2X2_6/Y gnd BUFX4_50/Y vdd BUFX4
XBUFX4_61 BUFX4_61/A gnd BUFX4_61/Y vdd BUFX4
XBUFX4_94 INVX8_1/Y gnd BUFX4_94/Y vdd BUFX4
XBUFX4_83 BUFX4_85/A gnd INVX8_13/A vdd BUFX4
XBUFX4_72 BUFX4_76/A gnd BUFX4_72/Y vdd BUFX4
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 INVX4_2/A INVX4_4/A gnd XNOR2X1_4/Y vdd XNOR2X1
XINVX8_20 INVX8_20/A gnd INVX8_20/Y vdd INVX8
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOAI21X1_562 BUFX4_148/Y OAI21X1_562/B BUFX4_164/Y gnd OAI22X1_115/D vdd OAI21X1
XOAI21X1_584 INVX4_10/A INVX8_22/Y INVX1_150/A gnd NOR2X1_231/B vdd OAI21X1
XOAI21X1_551 BUFX4_147/Y OAI21X1_551/B BUFX4_162/Y gnd OAI22X1_112/D vdd OAI21X1
XOAI21X1_540 INVX2_122/Y BUFX4_190/Y OAI21X1_617/C gnd OAI21X1_540/Y vdd OAI21X1
XOAI21X1_573 INVX2_65/Y MUX2X1_41/S OAI21X1_573/C gnd OAI21X1_573/Y vdd OAI21X1
XOAI21X1_595 BUFX4_121/Y INVX8_20/Y MUX2X1_24/Y gnd OAI21X1_596/C vdd OAI21X1
XFILL_22_0_1 gnd vdd FILL
XBUFX4_209 INVX8_8/Y gnd DFFSR_9/R vdd BUFX4
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_392 MUX2X1_8/A BUFX4_20/Y OAI21X1_641/C gnd OAI21X1_392/Y vdd OAI21X1
XOAI21X1_370 BUFX4_158/Y OAI21X1_370/B OAI21X1_370/C gnd AOI22X1_46/C vdd OAI21X1
XOAI21X1_381 OAI21X1_381/A BUFX4_244/Y OAI21X1_381/C gnd DFFSR_226/D vdd OAI21X1
XMUX2X1_16 MUX2X1_34/B MUX2X1_22/B MUX2X1_6/S gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_27 wb_dat_i[24] MUX2X1_27/B BUFX4_89/Y gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B MUX2X1_38/S gnd MUX2X1_38/Y vdd MUX2X1
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_9/R vdd DFFSR_8/D gnd vdd DFFSR
XNAND2X1_75 NOR2X1_38/Y NOR2X1_33/Y gnd OAI22X1_49/C vdd NAND2X1
XNAND2X1_86 INVX1_78/Y NOR3X1_1/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_20 BUFX4_25/Y wb_dat_i[11] gnd OAI21X1_99/C vdd NAND2X1
XNAND2X1_97 MUX2X1_2/Y NOR2X1_66/B gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_64 MUX2X1_19/B BUFX4_115/Y gnd NAND3X1_85/A vdd NAND2X1
XNAND2X1_53 INVX1_114/A BUFX4_116/Y gnd NAND3X1_74/A vdd NAND2X1
XNAND2X1_42 AOI21X1_8/Y NOR2X1_9/Y gnd DFFSR_72/D vdd NAND2X1
XNAND2X1_31 MUX2X1_35/S wb_dat_i[6] gnd OAI21X1_89/C vdd NAND2X1
XAOI21X1_224 NOR2X1_262/Y NOR2X1_259/B NOR2X1_263/Y gnd DFFSR_245/D vdd AOI21X1
XAOI21X1_202 INVX2_149/Y OAI21X1_579/B BUFX4_260/Y gnd OAI21X1_579/C vdd AOI21X1
XAOI21X1_213 NOR2X1_248/Y BUFX4_160/Y OAI21X1_680/Y gnd OAI22X1_120/C vdd AOI21X1
XAOI22X1_51 MUX2X1_4/A BUFX4_243/Y AOI22X1_51/C AOI22X1_51/D gnd DFFSR_223/D vdd AOI22X1
XAOI22X1_84 INVX2_69/Y BUFX4_5/Y AOI22X1_84/C AOI22X1_84/D gnd DFFSR_179/D vdd AOI22X1
XAOI22X1_62 INVX2_111/Y BUFX4_145/Y AOI22X1_62/C AOI22X1_62/D gnd DFFSR_202/D vdd
+ AOI22X1
XAOI22X1_73 INVX2_146/Y BUFX4_1/Y AOI22X1_73/C AOI22X1_73/D gnd DFFSR_164/D vdd AOI22X1
XAOI22X1_40 INVX2_115/Y BUFX4_246/Y AOI22X1_40/C AOI22X1_40/D gnd DFFSR_238/D vdd
+ AOI22X1
XNAND3X1_228 INVX2_140/Y BUFX4_49/Y BUFX4_138/Y gnd NAND3X1_229/C vdd NAND3X1
XNAND3X1_239 INVX2_145/Y BUFX4_71/Y BUFX4_61/Y gnd NAND3X1_241/B vdd NAND3X1
XNAND3X1_206 BUFX4_206/Y NAND3X1_206/B NAND3X1_206/C gnd AOI21X1_51/A vdd NAND3X1
XNAND3X1_217 BUFX4_204/Y NAND3X1_217/B NAND3X1_217/C gnd AOI21X1_52/A vdd NAND3X1
XOAI22X1_2 OAI22X1_5/A INVX2_10/Y INVX2_39/Y OAI22X1_5/D gnd NOR2X1_2/A vdd OAI22X1
XFILL_30_6_0 gnd vdd FILL
XDFFSR_248 INVX4_2/A CLKBUF1_41/Y BUFX4_15/Y vdd DFFSR_248/D gnd vdd DFFSR
XDFFSR_237 INVX2_84/A CLKBUF1_28/Y BUFX4_8/Y vdd DFFSR_237/D gnd vdd DFFSR
XDFFSR_204 INVX2_141/A CLKBUF1_40/Y BUFX4_17/Y vdd DFFSR_204/D gnd vdd DFFSR
XDFFSR_226 INVX2_106/A CLKBUF1_20/Y BUFX4_9/Y vdd DFFSR_226/D gnd vdd DFFSR
XDFFSR_215 INVX2_64/A CLKBUF1_1/Y BUFX4_16/Y vdd DFFSR_215/D gnd vdd DFFSR
XFILL_21_6_0 gnd vdd FILL
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XINVX2_44 INVX2_44/A gnd INVX2_44/Y vdd INVX2
XINVX2_11 DFFSR_2/Q gnd INVX2_11/Y vdd INVX2
XFILL_29_7_0 gnd vdd FILL
XINVX2_55 INVX2_55/A gnd INVX2_55/Y vdd INVX2
XINVX2_88 INVX2_88/A gnd INVX2_88/Y vdd INVX2
XINVX2_66 NOR3X1_4/B gnd INVX2_66/Y vdd INVX2
XFILL_4_7_0 gnd vdd FILL
XINVX2_99 INVX2_99/A gnd INVX2_99/Y vdd INVX2
XINVX2_77 INVX2_77/A gnd INVX2_77/Y vdd INVX2
XOAI21X1_29 INVX1_15/Y BUFX4_190/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XOAI21X1_18 BUFX4_102/Y INVX1_9/Y OAI21X1_18/C gnd DFFSR_17/D vdd OAI21X1
XFILL_12_6_0 gnd vdd FILL
XFILL_12_2 gnd vdd FILL
XNAND2X1_205 INVX8_17/A INVX1_145/Y gnd OAI21X1_410/B vdd NAND2X1
XNAND2X1_216 INVX4_12/A AND2X2_17/A gnd OAI21X1_547/B vdd NAND2X1
XNAND2X1_238 BUFX4_6/Y OAI21X1_641/Y gnd OAI21X1_643/C vdd NAND2X1
XNAND2X1_227 BUFX4_2/Y OAI21X1_609/Y gnd OAI21X1_612/C vdd NAND2X1
XNAND2X1_249 BUFX4_108/Y wb_dat_i[7] gnd OAI21X1_693/C vdd NAND2X1
XNOR2X1_260 NOR3X1_6/A INVX2_52/A gnd NOR2X1_260/Y vdd NOR2X1
XOAI21X1_711 NOR2X1_259/B OAI21X1_711/B OAI21X1_711/C gnd DFFSR_253/D vdd OAI21X1
XOAI21X1_700 OAI21X1_700/A BUFX4_1/Y OAI21X1_700/C gnd DFFSR_139/D vdd OAI21X1
XBUFX4_84 BUFX4_85/A gnd MUX2X1_9/S vdd BUFX4
XBUFX4_95 INVX8_1/Y gnd BUFX4_95/Y vdd BUFX4
XBUFX4_51 OR2X2_6/Y gnd BUFX4_51/Y vdd BUFX4
XBUFX4_73 BUFX4_76/A gnd BUFX4_73/Y vdd BUFX4
XBUFX4_62 BUFX4_66/A gnd BUFX4_62/Y vdd BUFX4
XCLKBUF1_19 CLKBUF1_6/A gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_40 BUFX4_45/A gnd INVX8_16/A vdd BUFX4
XOR2X2_10 OR2X2_10/A miso_pad_i gnd OR2X2_10/Y vdd OR2X2
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XXNOR2X1_5 XNOR2X1_5/A XOR2X1_2/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XINVX8_10 INVX8_10/A gnd INVX8_10/Y vdd INVX8
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XINVX8_21 BUFX4_2/Y gnd INVX8_21/Y vdd INVX8
XOAI21X1_530 AND2X2_19/Y INVX2_98/Y BUFX4_151/Y gnd OAI21X1_530/Y vdd OAI21X1
XOAI21X1_541 BUFX4_126/Y INVX2_156/Y INVX1_147/Y gnd NOR2X1_226/B vdd OAI21X1
XOAI21X1_552 NOR2X1_208/Y MUX2X1_15/A BUFX4_148/Y gnd OAI21X1_552/Y vdd OAI21X1
XOAI21X1_563 NOR2X1_211/Y INVX2_143/Y BUFX4_147/Y gnd OAI21X1_563/Y vdd OAI21X1
XOAI21X1_585 BUFX4_121/Y INVX8_20/Y MUX2X1_20/Y gnd OAI21X1_586/C vdd OAI21X1
XOAI21X1_574 BUFX4_159/Y OAI21X1_574/B OAI21X1_574/C gnd AOI22X1_80/C vdd OAI21X1
XOAI21X1_596 BUFX4_163/Y MUX2X1_23/Y OAI21X1_596/C gnd DFFSR_142/D vdd OAI21X1
.ends

