magic
tech scmos
timestamp 1751266522
<< metal1 >>
rect 896 3103 898 3107
rect 902 3103 905 3107
rect 909 3103 912 3107
rect 1928 3103 1930 3107
rect 1934 3103 1937 3107
rect 1941 3103 1944 3107
rect 2952 3103 2954 3107
rect 2958 3103 2961 3107
rect 2965 3103 2968 3107
rect 3976 3103 3978 3107
rect 3982 3103 3985 3107
rect 3989 3103 3992 3107
rect 618 3078 625 3081
rect 630 3071 633 3081
rect 3674 3078 3678 3082
rect 3766 3078 3777 3081
rect 630 3068 649 3071
rect 654 3068 665 3071
rect 806 3068 825 3071
rect 950 3071 953 3078
rect 3766 3072 3769 3078
rect 862 3068 873 3071
rect 910 3068 921 3071
rect 942 3068 953 3071
rect 1190 3068 1198 3071
rect 2070 3068 2086 3071
rect 3516 3068 3518 3072
rect 3790 3068 3801 3071
rect 654 3062 657 3068
rect 574 3058 593 3061
rect 910 3061 913 3068
rect 894 3058 913 3061
rect 1703 3058 1721 3061
rect 1975 3058 2009 3061
rect 3606 3058 3614 3061
rect 3670 3061 3673 3068
rect 3790 3062 3793 3068
rect 3638 3058 3673 3061
rect 3806 3061 3809 3071
rect 4038 3062 4041 3071
rect 3806 3058 3818 3061
rect 162 3048 169 3051
rect 574 3048 577 3058
rect 754 3048 756 3052
rect 954 3048 961 3051
rect 2606 3052 2610 3054
rect 3550 3051 3553 3058
rect 3814 3056 3818 3058
rect 3534 3048 3553 3051
rect 3718 3048 3729 3051
rect 3774 3046 3778 3048
rect 3486 3038 3502 3041
rect 3894 3041 3897 3061
rect 3930 3058 3937 3061
rect 3974 3058 3990 3061
rect 4058 3058 4065 3061
rect 4070 3058 4097 3061
rect 4222 3058 4230 3061
rect 4358 3058 4390 3061
rect 3982 3048 3990 3051
rect 3998 3048 4009 3051
rect 4046 3048 4057 3051
rect 3998 3042 4001 3048
rect 3894 3038 3921 3041
rect 4014 3038 4022 3041
rect 3605 3028 3606 3032
rect 826 3018 827 3022
rect 3637 3018 3638 3022
rect 3741 3018 3742 3022
rect 4154 3018 4155 3022
rect 392 3003 394 3007
rect 398 3003 401 3007
rect 405 3003 408 3007
rect 1416 3003 1418 3007
rect 1422 3003 1425 3007
rect 1429 3003 1432 3007
rect 2440 3003 2442 3007
rect 2446 3003 2449 3007
rect 2453 3003 2456 3007
rect 3472 3003 3474 3007
rect 3478 3003 3481 3007
rect 3485 3003 3488 3007
rect 2858 2988 2859 2992
rect 3165 2988 3166 2992
rect 3197 2988 3198 2992
rect 3997 2988 3998 2992
rect 1533 2978 1534 2982
rect 4110 2972 4113 2981
rect 374 2968 385 2971
rect 2573 2968 2574 2972
rect 2805 2968 2806 2972
rect 3570 2968 3571 2972
rect 3798 2968 3806 2971
rect 374 2966 378 2968
rect 374 2948 385 2951
rect 626 2948 641 2951
rect 646 2948 657 2951
rect 902 2948 937 2951
rect 990 2948 998 2951
rect 1418 2948 1449 2951
rect 1518 2951 1521 2961
rect 1502 2948 1521 2951
rect 2278 2951 2281 2961
rect 2262 2948 2281 2951
rect 2758 2951 2761 2958
rect 2758 2948 2769 2951
rect 374 2942 377 2948
rect 438 2941 441 2948
rect 654 2942 657 2948
rect 438 2938 457 2941
rect 550 2938 558 2941
rect 598 2938 606 2941
rect 978 2938 985 2941
rect 1010 2938 1017 2941
rect 1446 2938 1449 2948
rect 1970 2938 1985 2941
rect 2474 2938 2497 2941
rect 2790 2941 2793 2951
rect 2830 2948 2857 2951
rect 3150 2951 3153 2961
rect 3134 2948 3153 2951
rect 3398 2948 3409 2951
rect 3934 2948 3953 2951
rect 4022 2948 4030 2951
rect 4266 2948 4273 2951
rect 4330 2948 4337 2951
rect 4342 2948 4350 2951
rect 3406 2942 3409 2948
rect 2790 2938 2809 2941
rect 3782 2938 3801 2941
rect 3870 2938 3881 2941
rect 4318 2938 4329 2941
rect 622 2932 625 2938
rect 10 2928 17 2931
rect 370 2928 382 2931
rect 398 2928 414 2931
rect 558 2928 566 2931
rect 618 2928 625 2932
rect 1042 2928 1049 2931
rect 3414 2928 3422 2931
rect 3806 2928 3814 2931
rect 3838 2928 3846 2931
rect 3870 2931 3873 2938
rect 3862 2928 3873 2931
rect 3902 2928 3913 2931
rect 4150 2931 4153 2938
rect 4318 2932 4321 2938
rect 4142 2928 4153 2931
rect 570 2918 577 2921
rect 3532 2918 3534 2922
rect 4210 2918 4211 2922
rect 4229 2918 4230 2922
rect 896 2903 898 2907
rect 902 2903 905 2907
rect 909 2903 912 2907
rect 1928 2903 1930 2907
rect 1934 2903 1937 2907
rect 1941 2903 1944 2907
rect 2952 2903 2954 2907
rect 2958 2903 2961 2907
rect 2965 2903 2968 2907
rect 3976 2903 3978 2907
rect 3982 2903 3985 2907
rect 3989 2903 3992 2907
rect 874 2888 881 2891
rect 1010 2888 1012 2892
rect 1398 2888 1406 2891
rect 3586 2888 3587 2892
rect 3886 2888 3897 2891
rect 4170 2888 4172 2892
rect 3886 2882 3889 2888
rect 902 2878 918 2881
rect 1410 2878 1422 2881
rect 214 2868 225 2871
rect 598 2868 617 2871
rect 658 2868 673 2871
rect 1351 2868 1369 2871
rect 1830 2871 1833 2881
rect 2326 2878 2337 2881
rect 2334 2872 2337 2878
rect 3278 2872 3281 2881
rect 1814 2868 1833 2871
rect 2054 2868 2065 2871
rect 2294 2868 2305 2871
rect 2558 2868 2577 2871
rect 2590 2868 2601 2871
rect 2654 2868 2662 2871
rect 3254 2868 3265 2871
rect 3466 2868 3481 2871
rect 3542 2868 3550 2871
rect 3638 2868 3657 2871
rect 182 2858 201 2861
rect 262 2858 270 2861
rect 502 2861 505 2868
rect 502 2858 513 2861
rect 654 2858 662 2861
rect 894 2858 902 2861
rect 1070 2861 1073 2868
rect 1366 2862 1369 2868
rect 2590 2862 2593 2868
rect 1070 2858 1090 2861
rect 1546 2858 1553 2861
rect 2266 2858 2281 2861
rect 2646 2858 2654 2861
rect 2950 2861 2953 2868
rect 3262 2862 3265 2868
rect 2950 2858 2977 2861
rect 3246 2858 3254 2861
rect 3534 2858 3542 2861
rect 3602 2858 3609 2861
rect 3614 2858 3622 2861
rect 3686 2861 3689 2871
rect 3766 2871 3769 2878
rect 3758 2868 3769 2871
rect 3942 2862 3945 2871
rect 4118 2868 4126 2871
rect 4146 2868 4153 2871
rect 4274 2868 4289 2871
rect 4338 2868 4345 2871
rect 3686 2858 3705 2861
rect 3770 2858 3777 2861
rect 4014 2861 4017 2868
rect 4014 2858 4025 2861
rect 4078 2858 4097 2861
rect 4302 2858 4318 2861
rect 4326 2858 4350 2861
rect 4358 2858 4382 2861
rect 550 2848 569 2851
rect 862 2848 870 2851
rect 1398 2848 1406 2851
rect 3986 2848 3993 2851
rect 4034 2848 4041 2851
rect 4094 2848 4097 2858
rect 858 2838 881 2841
rect 1654 2838 1662 2841
rect 3666 2838 3667 2842
rect 4042 2838 4057 2841
rect 1846 2828 1854 2831
rect 13 2818 14 2822
rect 482 2818 483 2822
rect 589 2818 590 2822
rect 3740 2818 3742 2822
rect 392 2803 394 2807
rect 398 2803 401 2807
rect 405 2803 408 2807
rect 1416 2803 1418 2807
rect 1422 2803 1425 2807
rect 1429 2803 1432 2807
rect 2440 2803 2442 2807
rect 2446 2803 2449 2807
rect 2453 2803 2456 2807
rect 3472 2803 3474 2807
rect 3478 2803 3481 2807
rect 3485 2803 3488 2807
rect 586 2788 587 2792
rect 741 2788 742 2792
rect 2610 2788 2611 2792
rect 2653 2788 2654 2792
rect 2770 2788 2771 2792
rect 3506 2788 3507 2792
rect 538 2768 539 2772
rect 918 2768 937 2771
rect 1430 2768 1446 2771
rect 3098 2768 3099 2772
rect 3790 2768 3798 2771
rect 4110 2768 4121 2771
rect 18 2758 22 2762
rect 478 2758 486 2761
rect 918 2761 921 2768
rect 4110 2762 4113 2768
rect 22 2748 30 2751
rect 214 2748 233 2751
rect 322 2748 337 2751
rect 530 2748 537 2751
rect 578 2748 585 2751
rect 782 2751 785 2761
rect 910 2758 921 2761
rect 910 2752 913 2758
rect 766 2748 785 2751
rect 870 2748 881 2751
rect 922 2748 937 2751
rect 1022 2748 1033 2751
rect 1670 2748 1673 2758
rect 2578 2758 2582 2762
rect 3518 2758 3537 2761
rect 3678 2758 3686 2761
rect 4030 2758 4038 2761
rect 2154 2748 2161 2751
rect 2190 2748 2217 2751
rect 2518 2748 2534 2751
rect 2614 2748 2633 2751
rect 2690 2748 2697 2751
rect 2754 2748 2769 2751
rect 2826 2748 2833 2751
rect 3090 2748 3097 2751
rect 3798 2751 3801 2758
rect 3798 2748 3809 2751
rect 3842 2748 3849 2751
rect 3866 2748 3873 2751
rect 3918 2748 3929 2751
rect 4054 2751 4057 2761
rect 4130 2758 4137 2761
rect 3994 2748 4017 2751
rect 4054 2748 4073 2751
rect 4142 2748 4162 2751
rect 870 2742 873 2748
rect 1022 2742 1025 2748
rect 86 2738 94 2741
rect 166 2738 174 2741
rect 206 2738 217 2741
rect 246 2738 254 2741
rect 302 2738 310 2741
rect 506 2738 513 2741
rect 694 2738 713 2741
rect 1058 2738 1073 2741
rect 2190 2738 2198 2741
rect 2422 2738 2449 2741
rect 2678 2738 2694 2741
rect 2822 2738 2830 2741
rect 3319 2738 3337 2741
rect 3414 2738 3433 2741
rect 3558 2738 3574 2741
rect 3594 2738 3601 2741
rect 3742 2741 3745 2748
rect 3678 2738 3689 2741
rect 3726 2738 3745 2741
rect 3822 2738 3830 2741
rect 3862 2738 3870 2741
rect 3890 2738 3897 2741
rect 3926 2738 3929 2748
rect 4158 2746 4162 2748
rect 3950 2738 3969 2741
rect 4030 2738 4041 2741
rect 4066 2738 4073 2741
rect 4110 2738 4121 2741
rect 4222 2738 4225 2748
rect 4254 2741 4257 2751
rect 4250 2738 4257 2741
rect 102 2731 105 2738
rect 782 2732 785 2738
rect 102 2728 113 2731
rect 254 2728 265 2731
rect 782 2728 790 2732
rect 2854 2728 2865 2731
rect 3414 2728 3417 2738
rect 3758 2731 3761 2738
rect 3758 2728 3769 2731
rect 3874 2728 3881 2731
rect 3886 2728 3889 2738
rect 4258 2728 4265 2731
rect 2422 2718 2430 2721
rect 3364 2718 3366 2722
rect 3628 2718 3630 2722
rect 4354 2718 4356 2722
rect 896 2703 898 2707
rect 902 2703 905 2707
rect 909 2703 912 2707
rect 1928 2703 1930 2707
rect 1934 2703 1937 2707
rect 1941 2703 1944 2707
rect 2952 2703 2954 2707
rect 2958 2703 2961 2707
rect 2965 2703 2968 2707
rect 3976 2703 3978 2707
rect 3982 2703 3985 2707
rect 3989 2703 3992 2707
rect 894 2688 902 2691
rect 3802 2688 3803 2692
rect 218 2678 222 2682
rect 318 2672 321 2681
rect 374 2678 385 2681
rect 610 2678 625 2681
rect 954 2678 961 2681
rect 2806 2678 2814 2681
rect 3198 2678 3209 2681
rect 190 2668 209 2671
rect 270 2668 289 2671
rect 476 2668 505 2671
rect 206 2658 209 2668
rect 250 2658 257 2661
rect 342 2661 345 2668
rect 310 2658 329 2661
rect 342 2658 353 2661
rect 374 2658 377 2668
rect 590 2662 593 2671
rect 814 2671 817 2678
rect 814 2668 825 2671
rect 1831 2668 1846 2671
rect 2166 2668 2177 2671
rect 2278 2668 2289 2671
rect 2774 2668 2785 2671
rect 2166 2662 2169 2668
rect 934 2658 950 2661
rect 1230 2658 1257 2661
rect 1870 2658 1878 2661
rect 2330 2658 2337 2661
rect 2414 2661 2417 2668
rect 3110 2662 3113 2671
rect 3266 2668 3273 2671
rect 3538 2668 3545 2671
rect 3614 2668 3625 2671
rect 3694 2668 3702 2671
rect 3854 2671 3857 2681
rect 3854 2668 3873 2671
rect 3614 2662 3617 2668
rect 2414 2658 2433 2661
rect 2710 2658 2718 2661
rect 3054 2658 3062 2661
rect 3522 2658 3542 2661
rect 3546 2658 3553 2661
rect 3630 2658 3638 2661
rect 3702 2658 3710 2661
rect 3718 2658 3737 2661
rect 3886 2661 3889 2668
rect 3878 2658 3889 2661
rect 3934 2661 3937 2668
rect 4278 2662 4281 2671
rect 3926 2658 3937 2661
rect 4306 2658 4313 2661
rect 326 2648 329 2658
rect 906 2648 921 2651
rect 3734 2648 3737 2658
rect 1830 2638 1838 2641
rect 1954 2638 1969 2641
rect 3510 2638 3518 2641
rect 514 2618 515 2622
rect 3325 2618 3326 2622
rect 3898 2618 3899 2622
rect 4076 2618 4078 2622
rect 4362 2618 4364 2622
rect 392 2603 394 2607
rect 398 2603 401 2607
rect 405 2603 408 2607
rect 1416 2603 1418 2607
rect 1422 2603 1425 2607
rect 1429 2603 1432 2607
rect 2440 2603 2442 2607
rect 2446 2603 2449 2607
rect 2453 2603 2456 2607
rect 3472 2603 3474 2607
rect 3478 2603 3481 2607
rect 3485 2603 3488 2607
rect 821 2588 822 2592
rect 853 2588 854 2592
rect 2146 2588 2147 2592
rect 2274 2588 2275 2592
rect 2322 2588 2323 2592
rect 2522 2588 2523 2592
rect 2669 2588 2670 2592
rect 3114 2588 3115 2592
rect 3237 2588 3238 2592
rect 3954 2588 3955 2592
rect 590 2568 602 2571
rect 1798 2568 1806 2571
rect 598 2566 602 2568
rect 1798 2566 1802 2568
rect 1822 2566 1826 2568
rect 1518 2552 1521 2561
rect 2090 2558 2094 2562
rect 3266 2558 3270 2562
rect 3722 2558 3729 2561
rect 62 2548 89 2551
rect 118 2548 137 2551
rect 854 2548 862 2551
rect 1070 2548 1089 2551
rect 1118 2548 1126 2551
rect 86 2538 89 2548
rect 1430 2542 1433 2551
rect 1550 2551 1554 2554
rect 1550 2548 1569 2551
rect 150 2538 158 2541
rect 214 2538 225 2541
rect 614 2538 633 2541
rect 730 2538 737 2541
rect 862 2538 870 2541
rect 1126 2538 1145 2541
rect 1910 2538 1918 2541
rect 1974 2541 1977 2551
rect 2170 2548 2177 2551
rect 2206 2548 2225 2551
rect 2230 2548 2238 2551
rect 2362 2548 2377 2551
rect 2442 2548 2465 2551
rect 2494 2548 2505 2551
rect 2514 2548 2521 2551
rect 2630 2548 2641 2551
rect 2502 2542 2505 2548
rect 1958 2538 1977 2541
rect 2606 2541 2609 2548
rect 2910 2542 2913 2551
rect 3094 2548 3113 2551
rect 3310 2551 3313 2558
rect 3282 2548 3297 2551
rect 3310 2548 3329 2551
rect 3638 2548 3649 2551
rect 3782 2551 3785 2561
rect 4054 2561 4057 2568
rect 4046 2558 4057 2561
rect 3782 2548 3801 2551
rect 2606 2538 2625 2541
rect 2678 2538 2686 2541
rect 3094 2541 3097 2548
rect 3086 2538 3097 2541
rect 3158 2541 3161 2548
rect 3158 2538 3177 2541
rect 3222 2538 3230 2541
rect 3590 2538 3614 2541
rect 3642 2538 3649 2541
rect 3854 2541 3857 2551
rect 3970 2548 3993 2551
rect 4166 2551 4169 2561
rect 4130 2548 4145 2551
rect 4150 2548 4169 2551
rect 4182 2548 4209 2551
rect 3842 2538 3849 2541
rect 3854 2538 3865 2541
rect 3918 2538 3929 2541
rect 4366 2538 4374 2541
rect 214 2532 217 2538
rect 3862 2532 3865 2538
rect 158 2528 169 2531
rect 1046 2528 1065 2531
rect 1470 2528 1486 2531
rect 1978 2528 1985 2531
rect 2021 2528 2022 2532
rect 2574 2528 2585 2531
rect 2866 2528 2873 2531
rect 1794 2518 1795 2522
rect 1818 2518 1819 2522
rect 2293 2518 2294 2522
rect 4205 2518 4206 2522
rect 4300 2518 4302 2522
rect 4357 2518 4358 2522
rect 896 2503 898 2507
rect 902 2503 905 2507
rect 909 2503 912 2507
rect 1928 2503 1930 2507
rect 1934 2503 1937 2507
rect 1941 2503 1944 2507
rect 2952 2503 2954 2507
rect 2958 2503 2961 2507
rect 2965 2503 2968 2507
rect 3976 2503 3978 2507
rect 3982 2503 3985 2507
rect 3989 2503 3992 2507
rect 2365 2488 2366 2492
rect 3890 2488 3892 2492
rect 4189 2488 4190 2492
rect 166 2478 185 2481
rect 502 2478 510 2482
rect 3166 2478 3177 2481
rect 3458 2478 3473 2481
rect 3706 2478 3713 2481
rect 3790 2478 3801 2481
rect 4310 2478 4326 2481
rect 502 2472 505 2478
rect 3166 2472 3169 2478
rect 518 2468 529 2471
rect 1011 2468 1025 2471
rect 1410 2468 1433 2471
rect 1790 2468 1798 2471
rect 1834 2468 1841 2471
rect 2134 2468 2153 2471
rect 2262 2468 2273 2471
rect 2798 2468 2806 2471
rect 3042 2468 3057 2471
rect 1430 2462 1433 2468
rect 2262 2462 2265 2468
rect 198 2458 217 2461
rect 410 2458 417 2461
rect 598 2458 609 2461
rect 1242 2458 1249 2461
rect 1354 2458 1361 2461
rect 1590 2458 1609 2461
rect 1886 2458 1894 2461
rect 1922 2458 1950 2461
rect 1958 2458 1966 2461
rect 2206 2458 2214 2461
rect 2270 2458 2289 2461
rect 2766 2458 2774 2461
rect 3110 2461 3113 2468
rect 3366 2462 3369 2471
rect 3378 2468 3385 2471
rect 3494 2468 3513 2471
rect 3686 2468 3694 2471
rect 3714 2468 3721 2471
rect 3822 2468 3833 2471
rect 3986 2468 4001 2471
rect 4294 2468 4305 2471
rect 3494 2462 3497 2468
rect 3102 2458 3113 2461
rect 3218 2458 3233 2461
rect 3418 2458 3425 2461
rect 4082 2458 4089 2461
rect 4230 2461 4233 2468
rect 4230 2458 4249 2461
rect 4262 2458 4281 2461
rect 4350 2458 4358 2461
rect 606 2452 609 2458
rect 1590 2456 1594 2458
rect 1294 2448 1305 2451
rect 3202 2448 3206 2452
rect 4262 2448 4265 2458
rect 4162 2438 4163 2442
rect 2301 2418 2302 2422
rect 3900 2418 3902 2422
rect 4221 2418 4222 2422
rect 4250 2418 4251 2422
rect 392 2403 394 2407
rect 398 2403 401 2407
rect 405 2403 408 2407
rect 1416 2403 1418 2407
rect 1422 2403 1425 2407
rect 1429 2403 1432 2407
rect 2440 2403 2442 2407
rect 2446 2403 2449 2407
rect 2453 2403 2456 2407
rect 3472 2403 3474 2407
rect 3478 2403 3481 2407
rect 3485 2403 3488 2407
rect 1058 2388 1059 2392
rect 2858 2388 2859 2392
rect 2933 2388 2934 2392
rect 1125 2368 1126 2372
rect 1414 2368 1438 2371
rect 1658 2368 1659 2372
rect 2594 2368 2601 2371
rect 2642 2368 2643 2372
rect 3181 2368 3182 2372
rect 1414 2366 1418 2368
rect 1454 2366 1458 2368
rect 26 2348 41 2351
rect 726 2342 729 2351
rect 878 2348 881 2358
rect 1070 2358 1081 2361
rect 1362 2358 1369 2361
rect 1686 2358 1694 2361
rect 1750 2358 1761 2361
rect 1774 2358 1782 2361
rect 1750 2352 1753 2358
rect 1534 2348 1542 2351
rect 1638 2348 1646 2351
rect 1966 2348 1974 2351
rect 2062 2348 2070 2351
rect 2118 2348 2134 2351
rect 2462 2348 2470 2351
rect 2494 2351 2497 2361
rect 2494 2348 2513 2351
rect 2558 2351 2561 2361
rect 3326 2358 3337 2361
rect 2558 2348 2577 2351
rect 2902 2351 2905 2358
rect 3554 2358 3561 2361
rect 3570 2358 3574 2362
rect 3886 2358 3894 2361
rect 2902 2348 2921 2351
rect 3058 2348 3065 2351
rect 3842 2348 3849 2351
rect 4094 2351 4097 2361
rect 4186 2358 4190 2362
rect 4062 2348 4081 2351
rect 4094 2348 4113 2351
rect 4230 2351 4233 2361
rect 4230 2348 4249 2351
rect 14 2338 22 2341
rect 647 2338 665 2341
rect 1138 2338 1145 2341
rect 1914 2338 1945 2341
rect 1958 2338 1966 2341
rect 2034 2338 2041 2341
rect 2054 2338 2062 2341
rect 2094 2338 2102 2341
rect 2158 2338 2169 2341
rect 2198 2338 2217 2341
rect 2526 2338 2529 2348
rect 2622 2338 2630 2341
rect 2790 2338 2793 2348
rect 2806 2338 2817 2341
rect 2838 2338 2841 2348
rect 2942 2338 2977 2341
rect 3022 2341 3025 2348
rect 3022 2338 3041 2341
rect 3118 2338 3126 2341
rect 3254 2338 3270 2341
rect 3330 2338 3337 2341
rect 3974 2338 4009 2341
rect 4018 2338 4033 2341
rect 4078 2338 4081 2348
rect 4122 2338 4129 2341
rect 4166 2338 4177 2341
rect 4326 2338 4334 2341
rect 4362 2338 4369 2341
rect 22 2328 41 2331
rect 1766 2328 1769 2338
rect 3254 2328 3257 2338
rect 3282 2328 3286 2332
rect 4358 2328 4361 2338
rect 1410 2318 1411 2322
rect 1450 2318 1451 2322
rect 3834 2318 3835 2322
rect 3956 2318 3958 2322
rect 4090 2318 4091 2322
rect 896 2303 898 2307
rect 902 2303 905 2307
rect 909 2303 912 2307
rect 1928 2303 1930 2307
rect 1934 2303 1937 2307
rect 1941 2303 1944 2307
rect 2952 2303 2954 2307
rect 2958 2303 2961 2307
rect 2965 2303 2968 2307
rect 3976 2303 3978 2307
rect 3982 2303 3985 2307
rect 3989 2303 3992 2307
rect 1581 2288 1582 2292
rect 2438 2288 2454 2291
rect 3690 2288 3691 2292
rect 2382 2278 2390 2281
rect 4010 2278 4017 2281
rect 4298 2278 4305 2281
rect 626 2268 633 2271
rect 930 2268 937 2271
rect 1730 2268 1737 2271
rect 1798 2268 1814 2271
rect 1922 2268 1937 2271
rect 1994 2268 2001 2271
rect 2042 2268 2049 2271
rect 2342 2268 2361 2271
rect 2458 2268 2465 2271
rect 2554 2268 2561 2271
rect 3286 2268 3297 2271
rect 3382 2268 3390 2271
rect 3558 2268 3566 2271
rect 3682 2268 3689 2271
rect 3790 2268 3809 2271
rect 3998 2268 4014 2271
rect 4034 2268 4041 2271
rect 4198 2271 4201 2278
rect 4198 2268 4209 2271
rect 4226 2268 4233 2271
rect 4334 2268 4342 2271
rect 22 2258 34 2261
rect 78 2258 97 2261
rect 22 2252 25 2258
rect 30 2256 34 2258
rect 38 2248 50 2251
rect 462 2252 465 2262
rect 638 2258 657 2261
rect 674 2258 689 2261
rect 718 2258 726 2261
rect 838 2258 846 2261
rect 966 2258 993 2261
rect 1654 2258 1662 2261
rect 1830 2258 1838 2261
rect 1902 2258 1926 2261
rect 1958 2258 1966 2261
rect 2026 2258 2033 2261
rect 2110 2258 2126 2261
rect 2338 2258 2345 2261
rect 2398 2258 2406 2261
rect 2478 2258 2505 2261
rect 2570 2258 2577 2261
rect 2886 2258 2889 2268
rect 3078 2258 3081 2268
rect 3294 2262 3297 2268
rect 3254 2258 3262 2261
rect 3278 2258 3286 2261
rect 3530 2258 3553 2261
rect 3562 2258 3577 2261
rect 3674 2258 3681 2261
rect 3746 2258 3753 2261
rect 3822 2261 3825 2268
rect 3814 2258 3825 2261
rect 3870 2258 3890 2261
rect 4018 2258 4025 2261
rect 4274 2258 4281 2261
rect 3886 2256 3890 2258
rect 1346 2248 1353 2251
rect 2506 2248 2510 2252
rect 2518 2248 2537 2251
rect 2542 2248 2550 2251
rect 3422 2248 3433 2251
rect 3502 2248 3513 2251
rect 3562 2248 3569 2251
rect 3586 2248 3593 2251
rect 3658 2248 3662 2252
rect 4262 2248 4273 2251
rect 38 2242 41 2248
rect 46 2246 50 2248
rect 1038 2241 1042 2244
rect 870 2238 890 2241
rect 1030 2238 1042 2241
rect 1334 2238 1366 2241
rect 1574 2241 1578 2244
rect 1566 2238 1578 2241
rect 1682 2238 1683 2242
rect 1957 2238 1958 2242
rect 3525 2238 3526 2242
rect 4124 2238 4126 2242
rect 870 2228 873 2238
rect 3445 2228 3446 2232
rect 1845 2218 1846 2222
rect 2058 2218 2059 2222
rect 2085 2218 2086 2222
rect 3277 2218 3278 2222
rect 3954 2218 3955 2222
rect 4050 2218 4051 2222
rect 392 2203 394 2207
rect 398 2203 401 2207
rect 405 2203 408 2207
rect 1416 2203 1418 2207
rect 1422 2203 1425 2207
rect 1429 2203 1432 2207
rect 2440 2203 2442 2207
rect 2446 2203 2449 2207
rect 2453 2203 2456 2207
rect 3472 2203 3474 2207
rect 3478 2203 3481 2207
rect 3485 2203 3488 2207
rect 778 2188 779 2192
rect 1018 2188 1019 2192
rect 1069 2188 1070 2192
rect 3426 2188 3427 2192
rect 866 2168 878 2171
rect 954 2168 955 2172
rect 1358 2171 1361 2181
rect 4154 2178 4155 2182
rect 1342 2168 1361 2171
rect 4202 2168 4209 2171
rect 2094 2166 2098 2168
rect 3438 2158 3449 2161
rect 4226 2158 4230 2162
rect 270 2148 294 2151
rect 302 2148 310 2151
rect 326 2148 334 2151
rect 1322 2148 1329 2151
rect 1402 2148 1409 2151
rect 1734 2148 1742 2151
rect 1858 2148 1862 2151
rect 1974 2148 1982 2151
rect 2030 2148 2038 2151
rect 2178 2148 2185 2151
rect 2330 2148 2337 2151
rect 2498 2148 2513 2151
rect 2518 2148 2545 2151
rect 2550 2148 2558 2151
rect 2622 2148 2665 2151
rect 3166 2148 3177 2151
rect 3182 2148 3190 2151
rect 278 2138 286 2141
rect 1118 2141 1121 2148
rect 1090 2138 1097 2141
rect 1118 2138 1129 2141
rect 1134 2138 1142 2141
rect 1382 2138 1401 2141
rect 1666 2138 1673 2141
rect 1974 2138 1977 2148
rect 3166 2142 3169 2148
rect 2098 2138 2105 2141
rect 2134 2138 2145 2141
rect 2374 2138 2382 2141
rect 2458 2138 2481 2141
rect 2486 2138 2502 2141
rect 2622 2138 2630 2141
rect 2974 2138 2982 2141
rect 3186 2138 3193 2141
rect 3230 2138 3246 2141
rect 3302 2138 3318 2141
rect 3526 2138 3534 2141
rect 3750 2141 3753 2148
rect 4054 2142 4057 2151
rect 3742 2138 3753 2141
rect 3790 2138 3817 2141
rect 3834 2138 3849 2141
rect 3922 2138 3937 2141
rect 4330 2138 4337 2141
rect 510 2128 526 2131
rect 1606 2128 1614 2131
rect 1758 2131 1761 2138
rect 1750 2128 1761 2131
rect 3230 2128 3233 2138
rect 3302 2128 3305 2138
rect 3774 2132 3777 2138
rect 3886 2132 3889 2138
rect 3770 2128 3777 2132
rect 3882 2128 3889 2132
rect 3950 2128 3961 2131
rect 4182 2128 4201 2131
rect 4298 2118 4300 2122
rect 896 2103 898 2107
rect 902 2103 905 2107
rect 909 2103 912 2107
rect 1928 2103 1930 2107
rect 1934 2103 1937 2107
rect 1941 2103 1944 2107
rect 2952 2103 2954 2107
rect 2958 2103 2961 2107
rect 2965 2103 2968 2107
rect 3976 2103 3978 2107
rect 3982 2103 3985 2107
rect 3989 2103 3992 2107
rect 3490 2088 3497 2091
rect 3565 2088 3566 2092
rect 2114 2078 2121 2081
rect 3302 2078 3313 2081
rect 3906 2078 3918 2081
rect 62 2062 65 2071
rect 415 2068 446 2071
rect 1094 2068 1102 2071
rect 1614 2068 1622 2071
rect 1870 2062 1873 2071
rect 1910 2068 1918 2071
rect 1974 2068 1982 2071
rect 2038 2062 2041 2071
rect 2054 2068 2073 2071
rect 2102 2068 2110 2071
rect 2126 2068 2137 2071
rect 2406 2068 2417 2071
rect 2446 2068 2454 2071
rect 2954 2068 2969 2071
rect 2990 2068 3009 2071
rect 3338 2068 3353 2071
rect 3398 2068 3409 2071
rect 3670 2068 3681 2071
rect 3694 2068 3718 2071
rect 4038 2068 4065 2071
rect 4220 2068 4238 2071
rect 2126 2062 2129 2068
rect 3406 2062 3409 2068
rect 3678 2062 3681 2068
rect 22 2058 41 2061
rect 454 2058 470 2061
rect 478 2058 486 2061
rect 522 2058 529 2061
rect 946 2058 953 2061
rect 1010 2058 1017 2061
rect 1190 2058 1198 2061
rect 1410 2058 1433 2061
rect 1810 2058 1825 2061
rect 1982 2058 1990 2061
rect 2094 2058 2102 2061
rect 2486 2058 2513 2061
rect 2746 2058 2753 2061
rect 2802 2058 2809 2061
rect 2858 2058 2873 2061
rect 2918 2058 2926 2061
rect 2982 2058 2990 2061
rect 3230 2058 3246 2061
rect 3638 2058 3646 2061
rect 4330 2058 4337 2061
rect 4354 2058 4369 2061
rect 1166 2048 1177 2051
rect 2754 2048 2758 2052
rect 2810 2048 2814 2052
rect 2870 2048 2873 2058
rect 3230 2048 3233 2058
rect 3734 2048 3745 2051
rect 3754 2048 3758 2052
rect 4338 2048 4342 2052
rect 4350 2048 4353 2058
rect 742 2041 745 2048
rect 742 2038 753 2041
rect 1125 2038 1126 2042
rect 1029 2018 1030 2022
rect 1890 2018 1891 2022
rect 1949 2018 1950 2022
rect 4130 2018 4131 2022
rect 392 2003 394 2007
rect 398 2003 401 2007
rect 405 2003 408 2007
rect 1416 2003 1418 2007
rect 1422 2003 1425 2007
rect 1429 2003 1432 2007
rect 2440 2003 2442 2007
rect 2446 2003 2449 2007
rect 2453 2003 2456 2007
rect 3472 2003 3474 2007
rect 3478 2003 3481 2007
rect 3485 2003 3488 2007
rect 3661 1988 3662 1992
rect 3690 1988 3691 1992
rect 3714 1988 3715 1992
rect 642 1968 643 1972
rect 706 1968 742 1971
rect 930 1968 931 1972
rect 958 1971 961 1981
rect 942 1968 961 1971
rect 1134 1968 1146 1971
rect 1238 1971 1241 1981
rect 1162 1968 1185 1971
rect 1222 1968 1241 1971
rect 1306 1968 1307 1972
rect 4213 1968 4214 1972
rect 1142 1966 1146 1968
rect 1342 1966 1346 1968
rect 66 1958 70 1962
rect 98 1958 102 1962
rect 178 1958 182 1962
rect 718 1958 726 1961
rect 666 1948 673 1951
rect 678 1948 686 1951
rect 806 1948 814 1951
rect 894 1948 926 1951
rect 1278 1951 1281 1958
rect 1926 1958 1942 1961
rect 3106 1958 3110 1962
rect 3554 1958 3558 1962
rect 3566 1958 3577 1961
rect 1278 1948 1289 1951
rect 1374 1948 1382 1951
rect 1414 1948 1430 1951
rect 1682 1948 1689 1951
rect 1710 1948 1721 1951
rect 1938 1948 1953 1951
rect 2514 1948 2521 1951
rect 2526 1948 2553 1951
rect 230 1938 233 1948
rect 614 1938 617 1948
rect 982 1938 985 1948
rect 1718 1942 1721 1948
rect 2886 1942 2889 1951
rect 3018 1948 3041 1951
rect 3138 1948 3145 1951
rect 3502 1948 3510 1951
rect 3650 1948 3657 1951
rect 4014 1948 4033 1951
rect 4190 1948 4198 1951
rect 4294 1948 4305 1951
rect 4310 1948 4329 1951
rect 4014 1942 4017 1948
rect 4294 1942 4297 1948
rect 1146 1938 1153 1941
rect 1286 1938 1297 1941
rect 1762 1938 1769 1941
rect 2030 1938 2046 1941
rect 2466 1938 2473 1941
rect 3226 1938 3241 1941
rect 3458 1938 3489 1941
rect 3594 1938 3617 1941
rect 3682 1938 3689 1941
rect 3978 1938 4001 1941
rect 2082 1928 2089 1931
rect 2282 1928 2289 1931
rect 3454 1928 3457 1938
rect 3646 1928 3654 1931
rect 3670 1928 3678 1931
rect 4046 1928 4057 1931
rect 4074 1928 4081 1931
rect 1338 1918 1339 1922
rect 1725 1918 1726 1922
rect 1926 1918 1942 1921
rect 1989 1918 1990 1922
rect 4010 1918 4011 1922
rect 896 1903 898 1907
rect 902 1903 905 1907
rect 909 1903 912 1907
rect 1928 1903 1930 1907
rect 1934 1903 1937 1907
rect 1941 1903 1944 1907
rect 2952 1903 2954 1907
rect 2958 1903 2961 1907
rect 2965 1903 2968 1907
rect 3976 1903 3978 1907
rect 3982 1903 3985 1907
rect 3989 1903 3992 1907
rect 1605 1888 1606 1892
rect 2378 1888 2379 1892
rect 1754 1878 1761 1881
rect 3882 1878 3889 1881
rect 642 1868 649 1871
rect 838 1868 846 1871
rect 930 1868 937 1871
rect 1086 1868 1094 1871
rect 1690 1868 1697 1871
rect 1998 1868 2014 1871
rect 2066 1868 2073 1871
rect 2098 1868 2105 1871
rect 46 1858 54 1861
rect 70 1858 78 1861
rect 478 1852 481 1861
rect 714 1858 721 1861
rect 930 1858 945 1861
rect 1126 1858 1145 1861
rect 1226 1858 1233 1861
rect 1382 1858 1402 1861
rect 1962 1858 1985 1861
rect 2278 1861 2281 1871
rect 2334 1868 2353 1871
rect 2486 1868 2502 1871
rect 2738 1868 2753 1871
rect 3062 1868 3073 1871
rect 3122 1868 3129 1871
rect 3146 1868 3153 1871
rect 2334 1862 2337 1868
rect 2270 1858 2281 1861
rect 2314 1858 2321 1861
rect 2410 1858 2417 1861
rect 2422 1858 2438 1861
rect 3070 1861 3073 1868
rect 3182 1862 3185 1871
rect 3250 1868 3257 1871
rect 3070 1858 3086 1861
rect 3302 1861 3305 1871
rect 3562 1868 3569 1871
rect 3690 1868 3697 1871
rect 3826 1868 3849 1871
rect 3854 1868 3873 1871
rect 3990 1871 3994 1872
rect 3998 1871 4001 1878
rect 3990 1868 4001 1871
rect 4358 1868 4377 1871
rect 3302 1858 3329 1861
rect 3606 1858 3614 1861
rect 3670 1858 3678 1861
rect 3958 1858 3966 1861
rect 4062 1858 4070 1861
rect 4086 1861 4089 1868
rect 4086 1858 4097 1861
rect 1126 1856 1130 1858
rect 1398 1856 1402 1858
rect 670 1848 681 1851
rect 3326 1852 3329 1858
rect 3614 1848 3625 1851
rect 3798 1848 3809 1851
rect 278 1841 281 1848
rect 686 1846 690 1848
rect 270 1838 281 1841
rect 686 1838 694 1841
rect 786 1838 787 1842
rect 1110 1838 1126 1841
rect 1534 1841 1538 1844
rect 1526 1838 1538 1841
rect 1550 1841 1553 1848
rect 1598 1841 1602 1844
rect 1550 1838 1561 1841
rect 1590 1838 1602 1841
rect 4134 1838 4142 1841
rect 1018 1818 1019 1822
rect 1354 1818 1355 1822
rect 4058 1818 4059 1822
rect 392 1803 394 1807
rect 398 1803 401 1807
rect 405 1803 408 1807
rect 1416 1803 1418 1807
rect 1422 1803 1425 1807
rect 1429 1803 1432 1807
rect 2440 1803 2442 1807
rect 2446 1803 2449 1807
rect 2453 1803 2456 1807
rect 3472 1803 3474 1807
rect 3478 1803 3481 1807
rect 3485 1803 3488 1807
rect 1277 1788 1278 1792
rect 1658 1788 1659 1792
rect 2877 1788 2878 1792
rect 3261 1778 3262 1782
rect 1442 1768 1465 1771
rect 3362 1768 3363 1772
rect 4170 1768 4190 1771
rect 1230 1766 1234 1768
rect 434 1758 438 1762
rect 790 1758 798 1761
rect 1230 1758 1241 1761
rect 2074 1758 2078 1762
rect 2146 1758 2153 1761
rect 2270 1761 2273 1768
rect 2262 1758 2273 1761
rect 2474 1758 2478 1762
rect 2558 1758 2577 1761
rect 46 1748 65 1751
rect 1014 1748 1022 1751
rect 1086 1751 1090 1754
rect 1058 1748 1065 1751
rect 1070 1748 1090 1751
rect 1766 1748 1774 1751
rect 2090 1748 2105 1751
rect 2114 1748 2121 1751
rect 2194 1748 2201 1751
rect 2582 1751 2585 1761
rect 2826 1758 2830 1762
rect 2538 1748 2545 1751
rect 2582 1748 2601 1751
rect 791 1738 809 1741
rect 854 1738 862 1741
rect 942 1738 945 1748
rect 1174 1741 1177 1748
rect 2742 1742 2745 1751
rect 3166 1751 3169 1761
rect 3626 1758 3630 1762
rect 3166 1748 3182 1751
rect 3302 1751 3305 1758
rect 3302 1748 3321 1751
rect 3402 1748 3409 1751
rect 3434 1748 3449 1751
rect 3606 1748 3614 1751
rect 3670 1748 3686 1751
rect 1166 1738 1177 1741
rect 1694 1738 1702 1741
rect 2486 1738 2497 1741
rect 2518 1738 2537 1741
rect 2726 1738 2742 1741
rect 3110 1738 3121 1741
rect 3206 1738 3225 1741
rect 3270 1738 3273 1748
rect 3398 1738 3406 1741
rect 3510 1741 3513 1748
rect 3466 1738 3489 1741
rect 3510 1738 3521 1741
rect 3670 1738 3673 1748
rect 3786 1738 3801 1741
rect 3118 1732 3121 1738
rect 1970 1728 1977 1731
rect 2506 1728 2513 1731
rect 2678 1728 2689 1731
rect 3702 1728 3713 1731
rect 1245 1718 1246 1722
rect 2178 1718 2179 1722
rect 4158 1721 4161 1728
rect 4058 1718 4065 1721
rect 4150 1718 4161 1721
rect 896 1703 898 1707
rect 902 1703 905 1707
rect 909 1703 912 1707
rect 1928 1703 1930 1707
rect 1934 1703 1937 1707
rect 1941 1703 1944 1707
rect 2952 1703 2954 1707
rect 2958 1703 2961 1707
rect 2965 1703 2968 1707
rect 3976 1703 3978 1707
rect 3982 1703 3985 1707
rect 3989 1703 3992 1707
rect 2101 1688 2102 1692
rect 4020 1688 4022 1692
rect 506 1678 513 1681
rect 1442 1678 1449 1681
rect 1838 1672 1841 1681
rect 1854 1678 1862 1681
rect 2374 1678 2390 1681
rect 338 1668 345 1671
rect 402 1668 417 1671
rect 982 1668 993 1671
rect 1210 1668 1217 1671
rect 1374 1668 1385 1671
rect 1526 1668 1537 1671
rect 2022 1668 2030 1671
rect 2782 1668 2801 1671
rect 2854 1668 2865 1671
rect 3166 1668 3177 1671
rect 3210 1668 3217 1671
rect 3518 1671 3521 1681
rect 4070 1678 4081 1681
rect 4078 1672 4081 1678
rect 3470 1668 3505 1671
rect 3518 1668 3526 1671
rect 3562 1668 3569 1671
rect 3618 1668 3630 1671
rect 4226 1668 4233 1671
rect 4322 1668 4329 1671
rect 982 1662 985 1668
rect 1382 1662 1385 1668
rect 1534 1662 1537 1668
rect 46 1658 65 1661
rect 914 1658 929 1661
rect 954 1658 961 1661
rect 1198 1658 1206 1661
rect 1282 1658 1289 1661
rect 1326 1658 1334 1661
rect 1442 1658 1449 1661
rect 1642 1658 1649 1661
rect 1738 1658 1753 1661
rect 1870 1658 1897 1661
rect 1990 1658 2009 1661
rect 2062 1658 2065 1668
rect 2646 1658 2673 1661
rect 2754 1658 2761 1661
rect 3418 1658 3425 1661
rect 3558 1658 3566 1661
rect 4354 1658 4361 1661
rect 862 1648 873 1651
rect 1610 1648 1614 1652
rect 1810 1648 1814 1652
rect 1990 1648 1993 1658
rect 2166 1648 2174 1651
rect 2602 1648 2606 1652
rect 3578 1648 3582 1652
rect 3590 1648 3601 1651
rect 3722 1648 3726 1652
rect 4362 1648 4366 1652
rect 502 1641 505 1648
rect 1062 1642 1066 1644
rect 494 1638 505 1641
rect 702 1638 721 1641
rect 1126 1641 1130 1644
rect 1206 1641 1210 1644
rect 1334 1641 1338 1644
rect 1118 1638 1130 1641
rect 1198 1638 1210 1641
rect 1326 1638 1338 1641
rect 2178 1638 2185 1641
rect 3666 1638 3667 1642
rect 4006 1641 4009 1648
rect 3974 1638 4009 1641
rect 4202 1638 4209 1641
rect 4298 1638 4305 1641
rect 718 1628 721 1638
rect 392 1603 394 1607
rect 398 1603 401 1607
rect 405 1603 408 1607
rect 1416 1603 1418 1607
rect 1422 1603 1425 1607
rect 1429 1603 1432 1607
rect 2440 1603 2442 1607
rect 2446 1603 2449 1607
rect 2453 1603 2456 1607
rect 3472 1603 3474 1607
rect 3478 1603 3481 1607
rect 3485 1603 3488 1607
rect 698 1588 699 1592
rect 901 1588 902 1592
rect 1418 1588 1433 1591
rect 1570 1588 1571 1592
rect 1818 1588 1819 1592
rect 2170 1588 2171 1592
rect 3386 1588 3387 1592
rect 3501 1588 3502 1592
rect 130 1568 131 1572
rect 650 1568 651 1572
rect 1046 1568 1070 1571
rect 1158 1571 1161 1581
rect 3325 1578 3326 1582
rect 1142 1568 1161 1571
rect 1533 1568 1534 1572
rect 1602 1568 1603 1572
rect 1986 1568 1987 1572
rect 2194 1568 2201 1571
rect 2266 1568 2273 1571
rect 4050 1568 4062 1571
rect 4122 1568 4123 1572
rect 66 1558 70 1562
rect 806 1558 814 1561
rect 1298 1558 1302 1562
rect 1722 1558 1726 1562
rect 1766 1558 1774 1561
rect 46 1548 54 1551
rect 82 1548 89 1551
rect 642 1548 649 1551
rect 678 1548 694 1551
rect 786 1548 793 1551
rect 998 1548 1009 1551
rect 102 1538 121 1541
rect 402 1538 417 1541
rect 434 1538 441 1541
rect 634 1538 641 1541
rect 670 1538 673 1548
rect 1006 1542 1009 1548
rect 1254 1542 1257 1551
rect 1382 1548 1401 1551
rect 1502 1548 1510 1551
rect 1594 1548 1601 1551
rect 1726 1548 1734 1551
rect 1854 1548 1862 1551
rect 1918 1548 1950 1551
rect 1958 1548 1985 1551
rect 2026 1548 2033 1551
rect 2118 1548 2126 1551
rect 2142 1548 2169 1551
rect 2238 1551 2241 1561
rect 2222 1548 2241 1551
rect 2246 1548 2254 1551
rect 2310 1551 2313 1561
rect 2602 1558 2606 1562
rect 2294 1548 2313 1551
rect 2582 1548 2590 1551
rect 910 1538 918 1541
rect 922 1538 937 1541
rect 978 1538 985 1541
rect 1482 1538 1489 1541
rect 1666 1538 1673 1541
rect 1874 1538 1881 1541
rect 2654 1542 2657 1551
rect 2942 1548 2945 1558
rect 3626 1558 3630 1562
rect 3866 1558 3870 1562
rect 3878 1558 3889 1561
rect 3238 1548 3246 1551
rect 3326 1548 3334 1551
rect 3358 1548 3366 1551
rect 3514 1548 3521 1551
rect 3710 1548 3718 1551
rect 3850 1548 3865 1551
rect 3958 1548 3985 1551
rect 4070 1548 4081 1551
rect 4102 1548 4121 1551
rect 2198 1538 2209 1541
rect 2270 1538 2281 1541
rect 2326 1538 2334 1541
rect 2514 1538 2529 1541
rect 2670 1538 2686 1541
rect 2702 1538 2721 1541
rect 2766 1538 2782 1541
rect 3198 1538 3214 1541
rect 3442 1538 3449 1541
rect 3542 1538 3558 1541
rect 3638 1538 3649 1541
rect 3730 1538 3737 1541
rect 3742 1538 3761 1541
rect 3914 1538 3921 1541
rect 3998 1538 4006 1541
rect 4228 1538 4230 1542
rect 1406 1528 1414 1531
rect 3542 1528 3545 1538
rect 4158 1531 4161 1538
rect 4150 1528 4161 1531
rect 1098 1518 1105 1521
rect 2317 1518 2318 1522
rect 3470 1518 3478 1521
rect 896 1503 898 1507
rect 902 1503 905 1507
rect 909 1503 912 1507
rect 1928 1503 1930 1507
rect 1934 1503 1937 1507
rect 1941 1503 1944 1507
rect 2952 1503 2954 1507
rect 2958 1503 2961 1507
rect 2965 1503 2968 1507
rect 3976 1503 3978 1507
rect 3982 1503 3985 1507
rect 3989 1503 3992 1507
rect 853 1488 854 1492
rect 974 1488 982 1491
rect 1461 1488 1462 1492
rect 1506 1488 1507 1492
rect 1406 1478 1422 1481
rect 3782 1478 3793 1481
rect 4054 1478 4065 1481
rect 70 1468 81 1471
rect 474 1468 481 1471
rect 518 1468 526 1471
rect 878 1471 881 1478
rect 878 1468 892 1471
rect 914 1468 921 1471
rect 938 1468 945 1471
rect 1526 1468 1545 1471
rect 1774 1468 1793 1471
rect 1830 1471 1833 1478
rect 3790 1472 3793 1478
rect 4062 1472 4065 1478
rect 1830 1468 1841 1471
rect 1910 1468 1929 1471
rect 1990 1468 1998 1471
rect 2118 1468 2137 1471
rect 78 1462 81 1468
rect 2326 1462 2329 1471
rect 2338 1468 2345 1471
rect 2658 1468 2665 1471
rect 2678 1468 2686 1471
rect 3094 1468 3105 1471
rect 3114 1468 3129 1471
rect 3358 1462 3361 1471
rect 3450 1468 3465 1471
rect 3518 1468 3537 1471
rect 3610 1468 3617 1471
rect 3694 1468 3713 1471
rect 4132 1468 4153 1471
rect 4196 1468 4198 1472
rect 4254 1468 4273 1471
rect 22 1458 41 1461
rect 46 1458 54 1461
rect 58 1458 62 1461
rect 447 1458 478 1461
rect 498 1458 505 1461
rect 522 1458 537 1461
rect 658 1458 665 1461
rect 958 1458 969 1461
rect 1606 1458 1633 1461
rect 1702 1458 1729 1461
rect 1734 1458 1742 1461
rect 1862 1458 1889 1461
rect 2078 1458 2097 1461
rect 2110 1458 2118 1461
rect 2390 1458 2398 1461
rect 2686 1458 2694 1461
rect 2702 1458 2726 1461
rect 2746 1458 2753 1461
rect 3474 1458 3505 1461
rect 3606 1458 3609 1468
rect 3694 1462 3697 1468
rect 4166 1458 4169 1468
rect 870 1456 874 1458
rect 1410 1448 1433 1451
rect 2094 1448 2097 1458
rect 2106 1448 2110 1452
rect 2478 1451 2481 1458
rect 2470 1448 2481 1451
rect 3082 1448 3086 1452
rect 822 1442 826 1444
rect 1510 1442 1514 1444
rect 2021 1438 2022 1442
rect 538 1428 539 1432
rect 598 1428 601 1438
rect 730 1418 731 1422
rect 1749 1418 1750 1422
rect 2818 1418 2819 1422
rect 2842 1418 2843 1422
rect 2870 1418 2878 1421
rect 3733 1418 3734 1422
rect 392 1403 394 1407
rect 398 1403 401 1407
rect 405 1403 408 1407
rect 1416 1403 1418 1407
rect 1422 1403 1425 1407
rect 1429 1403 1432 1407
rect 2440 1403 2442 1407
rect 2446 1403 2449 1407
rect 2453 1403 2456 1407
rect 3472 1403 3474 1407
rect 3478 1403 3481 1407
rect 3485 1403 3488 1407
rect 770 1388 771 1392
rect 1210 1388 1211 1392
rect 1253 1388 1254 1392
rect 1906 1388 1907 1392
rect 2069 1388 2070 1392
rect 3405 1388 3406 1392
rect 4106 1388 4107 1392
rect 4330 1388 4331 1392
rect 798 1372 801 1381
rect 66 1368 67 1372
rect 866 1368 873 1371
rect 3834 1368 3835 1372
rect 686 1366 690 1368
rect 122 1358 126 1362
rect 898 1358 902 1362
rect 946 1358 950 1362
rect 1078 1358 1086 1361
rect 1434 1358 1441 1361
rect 58 1348 65 1351
rect 302 1348 305 1358
rect 494 1348 497 1358
rect 718 1348 734 1351
rect 826 1348 833 1351
rect 930 1348 945 1351
rect 1118 1348 1137 1351
rect 1190 1348 1209 1351
rect 1382 1348 1401 1351
rect 1622 1348 1649 1351
rect 1678 1348 1686 1351
rect 1710 1351 1713 1361
rect 1874 1358 1878 1362
rect 1918 1358 1926 1361
rect 2298 1358 2302 1362
rect 2442 1358 2457 1361
rect 2526 1358 2537 1361
rect 2682 1358 2686 1362
rect 2694 1358 2705 1361
rect 3330 1358 3334 1362
rect 3846 1358 3857 1361
rect 4126 1358 4129 1368
rect 1710 1348 1729 1351
rect 1754 1348 1761 1351
rect 1846 1351 1849 1358
rect 1830 1348 1849 1351
rect 2358 1348 2369 1351
rect 2558 1348 2566 1351
rect 2818 1348 2825 1351
rect 2934 1348 2966 1351
rect 2982 1348 3009 1351
rect 3254 1348 3262 1351
rect 3394 1348 3401 1351
rect 3742 1348 3753 1351
rect 3814 1348 3822 1351
rect 710 1338 713 1348
rect 1190 1341 1193 1348
rect 1182 1338 1193 1341
rect 1262 1338 1270 1341
rect 1382 1341 1385 1348
rect 1374 1338 1385 1341
rect 1502 1338 1521 1341
rect 1582 1338 1601 1341
rect 1782 1338 1801 1341
rect 1990 1341 1993 1348
rect 1930 1338 1953 1341
rect 1990 1338 2001 1341
rect 2390 1338 2417 1341
rect 2422 1338 2457 1341
rect 2530 1338 2537 1341
rect 2558 1338 2561 1348
rect 2590 1338 2609 1341
rect 2622 1338 2641 1341
rect 2722 1338 2745 1341
rect 2878 1341 2881 1348
rect 2870 1338 2881 1341
rect 2894 1338 2913 1341
rect 2954 1338 2969 1341
rect 3342 1338 3350 1341
rect 3390 1338 3398 1341
rect 3662 1338 3681 1341
rect 3814 1338 3817 1348
rect 4022 1342 4025 1351
rect 4270 1348 4278 1351
rect 4322 1348 4329 1351
rect 3972 1338 4009 1341
rect 4214 1338 4217 1348
rect 4366 1338 4374 1341
rect 682 1328 694 1331
rect 1142 1328 1145 1338
rect 2622 1332 2625 1338
rect 3662 1332 3665 1338
rect 2082 1328 2089 1331
rect 3414 1328 3422 1331
rect 3742 1328 3750 1331
rect 1314 1318 1315 1322
rect 4148 1318 4150 1322
rect 896 1303 898 1307
rect 902 1303 905 1307
rect 909 1303 912 1307
rect 1928 1303 1930 1307
rect 1934 1303 1937 1307
rect 1941 1303 1944 1307
rect 2952 1303 2954 1307
rect 2958 1303 2961 1307
rect 2965 1303 2968 1307
rect 3976 1303 3978 1307
rect 3982 1303 3985 1307
rect 3989 1303 3992 1307
rect 1085 1288 1086 1292
rect 1926 1288 1942 1291
rect 3956 1288 3966 1291
rect 1442 1278 1449 1281
rect 343 1268 358 1271
rect 774 1268 790 1271
rect 1422 1268 1446 1271
rect 1454 1268 1473 1271
rect 1566 1262 1569 1271
rect 1626 1268 1633 1271
rect 1686 1271 1689 1281
rect 1662 1268 1681 1271
rect 1686 1268 1702 1271
rect 1786 1268 1793 1271
rect 1938 1268 1961 1271
rect 2026 1268 2033 1271
rect 3022 1268 3033 1271
rect 3062 1268 3081 1271
rect 3094 1268 3105 1271
rect 3238 1268 3246 1271
rect 3270 1271 3273 1281
rect 3298 1278 3302 1282
rect 3382 1278 3390 1282
rect 3382 1272 3385 1278
rect 3270 1268 3286 1271
rect 3430 1271 3433 1281
rect 3430 1268 3446 1271
rect 3474 1268 3497 1271
rect 3550 1271 3553 1281
rect 3638 1278 3646 1281
rect 3924 1278 3926 1282
rect 4298 1278 4305 1281
rect 3550 1268 3569 1271
rect 4022 1271 4025 1278
rect 4022 1268 4036 1271
rect 4246 1271 4250 1272
rect 4254 1271 4257 1278
rect 4164 1268 4185 1271
rect 4246 1268 4257 1271
rect 3094 1262 3097 1268
rect 366 1258 385 1261
rect 598 1258 606 1261
rect 1494 1258 1502 1261
rect 1514 1258 1521 1261
rect 1622 1258 1630 1261
rect 1726 1258 1734 1261
rect 1870 1258 1889 1261
rect 1954 1258 1961 1261
rect 2006 1258 2014 1261
rect 2286 1258 2294 1261
rect 2734 1258 2742 1261
rect 3106 1258 3113 1261
rect 3166 1258 3174 1261
rect 3242 1258 3249 1261
rect 3470 1258 3478 1261
rect 3662 1258 3670 1261
rect 4070 1258 4081 1261
rect 398 1248 414 1251
rect 606 1248 614 1251
rect 710 1248 721 1251
rect 1490 1248 1494 1252
rect 1926 1248 1934 1251
rect 2062 1251 2065 1258
rect 2062 1248 2073 1251
rect 2754 1248 2758 1252
rect 2766 1248 2777 1251
rect 3114 1248 3118 1252
rect 3162 1248 3166 1252
rect 3330 1248 3334 1252
rect 3518 1248 3521 1258
rect 3718 1248 3729 1251
rect 3806 1248 3817 1251
rect 694 1242 698 1244
rect 666 1238 673 1241
rect 710 1242 713 1248
rect 966 1242 970 1244
rect 3382 1242 3386 1244
rect 726 1238 734 1241
rect 1162 1238 1169 1241
rect 3229 1228 3230 1232
rect 3506 1228 3507 1232
rect 813 1218 814 1222
rect 1298 1218 1299 1222
rect 1330 1218 1331 1222
rect 1586 1218 1587 1222
rect 3658 1218 3659 1222
rect 3706 1218 3707 1222
rect 3765 1218 3766 1222
rect 392 1203 394 1207
rect 398 1203 401 1207
rect 405 1203 408 1207
rect 1416 1203 1418 1207
rect 1422 1203 1425 1207
rect 1429 1203 1432 1207
rect 2440 1203 2442 1207
rect 2446 1203 2449 1207
rect 2453 1203 2456 1207
rect 3472 1203 3474 1207
rect 3478 1203 3481 1207
rect 3485 1203 3488 1207
rect 1506 1188 1507 1192
rect 1554 1188 1555 1192
rect 1618 1188 1619 1192
rect 1682 1188 1683 1192
rect 1909 1188 1910 1192
rect 3130 1188 3131 1192
rect 3378 1188 3379 1192
rect 3974 1188 3990 1191
rect 4138 1188 4139 1192
rect 390 1178 398 1181
rect 918 1172 921 1181
rect 4326 1172 4329 1181
rect 578 1168 593 1171
rect 650 1168 651 1172
rect 870 1166 874 1168
rect 866 1158 873 1161
rect 878 1158 913 1161
rect 1718 1158 1726 1161
rect 1978 1158 1982 1162
rect 2842 1158 2846 1162
rect 3034 1158 3038 1162
rect 3390 1158 3401 1161
rect 4278 1158 4294 1161
rect 26 1148 33 1151
rect 130 1148 137 1151
rect 374 1148 382 1151
rect 458 1148 473 1151
rect 962 1148 969 1151
rect 998 1148 1006 1151
rect 1134 1148 1142 1151
rect 1398 1148 1422 1151
rect 1486 1148 1494 1151
rect 1510 1148 1518 1151
rect 1654 1148 1670 1151
rect 1686 1148 1702 1151
rect 1958 1148 1966 1151
rect 1982 1148 1998 1151
rect 2886 1148 2913 1151
rect 3038 1148 3065 1151
rect 3746 1148 3753 1151
rect 3894 1148 3905 1151
rect 30 1138 33 1148
rect 4086 1142 4089 1151
rect 66 1138 73 1141
rect 110 1138 126 1141
rect 162 1138 169 1141
rect 454 1138 462 1141
rect 610 1138 617 1141
rect 734 1138 742 1141
rect 886 1138 902 1141
rect 1322 1138 1329 1141
rect 1458 1138 1465 1141
rect 1774 1138 1790 1141
rect 1862 1138 1870 1141
rect 1962 1138 1969 1141
rect 2574 1138 2593 1141
rect 2958 1138 2974 1141
rect 3138 1138 3150 1141
rect 3246 1138 3254 1141
rect 3258 1138 3262 1141
rect 3318 1138 3334 1141
rect 3918 1138 3937 1141
rect 1102 1132 1105 1138
rect 1098 1128 1105 1132
rect 2014 1131 2017 1138
rect 2006 1128 2017 1131
rect 3166 1128 3177 1131
rect 3246 1128 3249 1138
rect 3318 1128 3321 1138
rect 3474 1128 3486 1131
rect 896 1103 898 1107
rect 902 1103 905 1107
rect 909 1103 912 1107
rect 1928 1103 1930 1107
rect 1934 1103 1937 1107
rect 1941 1103 1944 1107
rect 2952 1103 2954 1107
rect 2958 1103 2961 1107
rect 2965 1103 2968 1107
rect 3976 1103 3978 1107
rect 3982 1103 3985 1107
rect 3989 1103 3992 1107
rect 3557 1088 3558 1092
rect 3717 1088 3718 1092
rect 4092 1088 4094 1092
rect 4206 1088 4217 1091
rect 4252 1088 4254 1092
rect 4206 1082 4209 1088
rect 986 1078 993 1081
rect 1406 1078 1422 1081
rect 2166 1078 2174 1081
rect 2970 1078 2977 1081
rect 3198 1078 3206 1081
rect 3482 1078 3489 1081
rect 3686 1078 3697 1081
rect 2534 1076 2538 1078
rect 615 1068 633 1071
rect 1026 1068 1033 1071
rect 1314 1068 1321 1071
rect 1462 1068 1470 1071
rect 46 1058 65 1061
rect 234 1058 241 1061
rect 246 1058 254 1061
rect 422 1052 425 1061
rect 638 1058 654 1061
rect 1478 1061 1481 1071
rect 1510 1068 1529 1071
rect 1966 1068 1985 1071
rect 1994 1068 2001 1071
rect 2126 1068 2134 1071
rect 3190 1068 3198 1071
rect 3226 1068 3233 1071
rect 3318 1068 3326 1071
rect 3410 1068 3417 1071
rect 3570 1068 3585 1071
rect 3590 1068 3617 1071
rect 3654 1068 3662 1071
rect 3678 1068 3689 1071
rect 3746 1068 3761 1071
rect 3948 1068 3950 1072
rect 3966 1071 3970 1072
rect 3974 1071 3977 1078
rect 3966 1068 3977 1071
rect 4142 1071 4146 1072
rect 4150 1071 4153 1078
rect 4142 1068 4153 1071
rect 4286 1068 4294 1071
rect 1474 1058 1481 1061
rect 1538 1058 1553 1061
rect 1658 1058 1665 1061
rect 1678 1058 1702 1061
rect 1786 1058 1793 1061
rect 1882 1058 1889 1061
rect 2402 1058 2409 1061
rect 2414 1058 2430 1061
rect 2442 1058 2449 1061
rect 2590 1058 2598 1061
rect 2878 1058 2886 1061
rect 2910 1058 2937 1061
rect 3210 1058 3217 1061
rect 3230 1058 3233 1068
rect 3310 1058 3334 1061
rect 3646 1061 3649 1068
rect 3686 1062 3689 1068
rect 3638 1058 3649 1061
rect 254 1048 273 1051
rect 658 1048 662 1052
rect 754 1048 758 1052
rect 1497 1048 1502 1052
rect 1586 1048 1590 1052
rect 1662 1048 1665 1058
rect 2086 1048 2105 1051
rect 2970 1048 2977 1051
rect 3370 1048 3374 1052
rect 3978 1038 4017 1041
rect 4014 1028 4017 1038
rect 1957 1018 1958 1022
rect 2858 1018 2859 1022
rect 392 1003 394 1007
rect 398 1003 401 1007
rect 405 1003 408 1007
rect 1416 1003 1418 1007
rect 1422 1003 1425 1007
rect 1429 1003 1432 1007
rect 2440 1003 2442 1007
rect 2446 1003 2449 1007
rect 2453 1003 2456 1007
rect 3472 1003 3474 1007
rect 3478 1003 3481 1007
rect 3485 1003 3488 1007
rect 1573 988 1574 992
rect 1629 988 1630 992
rect 1810 988 1811 992
rect 1901 988 1902 992
rect 1934 988 1942 991
rect 2690 988 2691 992
rect 4290 988 4291 992
rect 1994 978 1995 982
rect 2746 968 2753 971
rect 4250 968 4265 971
rect 1022 966 1026 968
rect 242 958 246 962
rect 1722 958 1729 961
rect 2626 958 2630 962
rect 2638 958 2649 961
rect 2702 958 2713 961
rect 2854 958 2862 961
rect 3594 958 3598 962
rect 3934 958 3945 961
rect 46 948 65 951
rect 278 948 286 951
rect 662 948 681 951
rect 906 948 929 951
rect 1070 942 1073 951
rect 1486 948 1494 951
rect 1630 948 1657 951
rect 1662 948 1670 951
rect 1702 948 1710 951
rect 1962 948 1969 951
rect 2006 948 2030 951
rect 2062 948 2070 951
rect 2450 948 2465 951
rect 2470 948 2478 951
rect 2890 948 2897 951
rect 3142 948 3161 951
rect 3522 948 3529 951
rect 3566 948 3590 951
rect 3926 948 3934 951
rect 4366 948 4374 951
rect 694 938 705 941
rect 954 938 961 941
rect 1034 938 1041 941
rect 1054 938 1062 941
rect 1234 938 1241 941
rect 1546 938 1553 941
rect 2026 938 2033 941
rect 2406 941 2409 948
rect 2406 938 2417 941
rect 2726 938 2734 941
rect 2826 938 2833 941
rect 2886 938 2889 948
rect 2910 938 2934 941
rect 3142 938 3145 948
rect 3182 938 3190 941
rect 3430 938 3438 941
rect 3442 938 3446 941
rect 3542 938 3550 941
rect 3662 938 3670 941
rect 3734 938 3742 941
rect 702 932 705 938
rect 1125 928 1126 932
rect 1378 928 1379 932
rect 1414 928 1430 931
rect 3430 928 3433 938
rect 1018 918 1019 922
rect 3389 918 3390 922
rect 3786 918 3787 922
rect 896 903 898 907
rect 902 903 905 907
rect 909 903 912 907
rect 1928 903 1930 907
rect 1934 903 1937 907
rect 1941 903 1944 907
rect 2952 903 2954 907
rect 2958 903 2961 907
rect 2965 903 2968 907
rect 3976 903 3978 907
rect 3982 903 3985 907
rect 3989 903 3992 907
rect 1234 888 1235 892
rect 1282 888 1283 892
rect 2438 888 2446 891
rect 2661 888 2662 892
rect 4046 888 4054 891
rect 4282 888 4284 892
rect 4346 888 4348 892
rect 1050 878 1057 881
rect 1434 878 1441 881
rect 2074 878 2081 881
rect 2122 878 2129 881
rect 2986 878 2993 881
rect 4118 881 4121 888
rect 4110 878 4121 881
rect 326 868 334 871
rect 1446 868 1454 871
rect 1470 868 1489 871
rect 1518 868 1529 871
rect 1670 868 1681 871
rect 1846 868 1857 871
rect 2554 868 2577 871
rect 2702 868 2710 871
rect 2714 868 2721 871
rect 3138 868 3145 871
rect 3278 868 3297 871
rect 3430 868 3438 871
rect 3738 868 3745 871
rect 3866 868 3889 871
rect 4092 868 4094 872
rect 4162 868 4177 871
rect 1670 862 1673 868
rect 1766 862 1770 864
rect 1846 862 1849 868
rect 690 858 705 861
rect 802 858 817 861
rect 1354 858 1361 861
rect 1578 858 1601 861
rect 1718 858 1745 861
rect 1810 858 1817 861
rect 2382 858 2401 861
rect 2702 858 2705 868
rect 2854 858 2870 861
rect 2886 858 2913 861
rect 2962 858 2990 861
rect 3006 858 3033 861
rect 3134 858 3142 861
rect 3178 858 3185 861
rect 3506 858 3513 861
rect 3830 858 3838 861
rect 1362 848 1366 852
rect 1618 848 1625 851
rect 2382 848 2385 858
rect 2526 848 2537 851
rect 2946 848 2951 852
rect 3330 848 3334 852
rect 3374 848 3385 851
rect 3838 848 3849 851
rect 3982 848 3998 851
rect 1238 842 1242 844
rect 242 838 243 842
rect 1286 842 1290 844
rect 1306 838 1307 842
rect 1602 838 1603 842
rect 2350 838 2358 841
rect 3974 838 4014 841
rect 3362 828 3363 832
rect 3974 828 3977 838
rect 1573 818 1574 822
rect 1637 818 1638 822
rect 2842 818 2843 822
rect 392 803 394 807
rect 398 803 401 807
rect 405 803 408 807
rect 1416 803 1418 807
rect 1422 803 1425 807
rect 1429 803 1432 807
rect 2440 803 2442 807
rect 2446 803 2449 807
rect 2453 803 2456 807
rect 3472 803 3474 807
rect 3478 803 3481 807
rect 3485 803 3488 807
rect 1434 788 1441 791
rect 1506 788 1507 792
rect 1538 788 1539 792
rect 1586 788 1587 792
rect 1674 788 1675 792
rect 1706 788 1707 792
rect 1738 788 1739 792
rect 1805 788 1806 792
rect 2050 788 2051 792
rect 314 768 315 772
rect 758 768 766 771
rect 2602 768 2609 771
rect 2653 768 2654 772
rect 3522 768 3523 772
rect 3830 768 3838 771
rect 686 758 697 761
rect 1174 761 1177 768
rect 1174 758 1185 761
rect 46 748 65 751
rect 626 748 633 751
rect 698 748 705 751
rect 710 748 718 751
rect 1522 748 1537 751
rect 1654 748 1662 751
rect 1750 751 1753 761
rect 2018 758 2022 762
rect 2590 758 2598 761
rect 2898 758 2902 762
rect 2946 758 2958 761
rect 3534 758 3545 761
rect 3894 758 3910 761
rect 3970 758 3985 761
rect 1750 748 1761 751
rect 1926 748 1934 751
rect 1970 748 1977 751
rect 2366 748 2377 751
rect 2430 748 2446 751
rect 2922 748 2929 751
rect 3254 748 3265 751
rect 726 738 729 748
rect 750 738 761 741
rect 1054 738 1073 741
rect 1146 738 1158 741
rect 1174 738 1177 748
rect 1758 741 1761 748
rect 1758 738 1769 741
rect 1930 738 1953 741
rect 2262 738 2270 741
rect 2662 738 2670 741
rect 2870 738 2878 741
rect 3030 738 3046 741
rect 3222 738 3233 741
rect 3222 732 3225 738
rect 3798 732 3801 738
rect 1414 728 1430 731
rect 1862 728 1870 731
rect 3794 728 3801 732
rect 1165 718 1166 722
rect 2397 718 2398 722
rect 3701 718 3702 722
rect 896 703 898 707
rect 902 703 905 707
rect 909 703 912 707
rect 1928 703 1930 707
rect 1934 703 1937 707
rect 1941 703 1944 707
rect 2952 703 2954 707
rect 2958 703 2961 707
rect 2965 703 2968 707
rect 3976 703 3978 707
rect 3982 703 3985 707
rect 3989 703 3992 707
rect 2645 688 2646 692
rect 3914 688 3921 691
rect 3990 688 3998 691
rect 4218 688 4225 691
rect 1750 678 1761 681
rect 2394 678 2409 681
rect 3362 678 3369 681
rect 3646 678 3657 681
rect 1750 672 1753 678
rect 790 668 801 671
rect 1574 668 1593 671
rect 2318 668 2329 671
rect 2606 668 2614 671
rect 2858 668 2865 671
rect 2886 668 2897 671
rect 2926 668 2937 671
rect 3534 668 3542 671
rect 3834 668 3841 671
rect 4126 671 4129 678
rect 4116 668 4129 671
rect 4170 668 4185 671
rect 4286 671 4290 672
rect 4282 668 4290 671
rect 4362 668 4377 671
rect 22 658 41 661
rect 890 658 913 661
rect 938 658 945 661
rect 1218 658 1225 661
rect 1326 658 1345 661
rect 1354 658 1369 661
rect 1394 658 1401 661
rect 1442 658 1462 661
rect 1542 658 1569 661
rect 1574 658 1577 668
rect 2318 662 2321 668
rect 2886 662 2889 668
rect 1638 658 1665 661
rect 2246 658 2273 661
rect 2290 658 2297 661
rect 2330 658 2337 661
rect 2374 658 2390 661
rect 2774 658 2798 661
rect 3506 658 3521 661
rect 3538 658 3545 661
rect 1326 656 1330 658
rect 2338 648 2342 652
rect 2802 648 2806 652
rect 3002 648 3006 652
rect 3402 648 3406 652
rect 3846 651 3849 658
rect 3846 648 3857 651
rect 3622 638 3630 641
rect 3646 641 3649 648
rect 3638 638 3649 641
rect 4002 638 4022 641
rect 4218 638 4225 641
rect 3810 628 3811 632
rect 3974 631 3977 638
rect 3958 628 3977 631
rect 4062 628 4065 638
rect 1786 618 1787 622
rect 1918 618 1934 621
rect 2621 618 2622 622
rect 2674 618 2675 622
rect 2709 618 2710 622
rect 3354 618 3355 622
rect 3378 618 3379 622
rect 392 603 394 607
rect 398 603 401 607
rect 405 603 408 607
rect 1416 603 1418 607
rect 1422 603 1425 607
rect 1429 603 1432 607
rect 2440 603 2442 607
rect 2446 603 2449 607
rect 2453 603 2456 607
rect 3472 603 3474 607
rect 3478 603 3481 607
rect 3485 603 3488 607
rect 1461 588 1462 592
rect 1490 588 1491 592
rect 1522 588 1523 592
rect 1650 588 1651 592
rect 1725 588 1726 592
rect 1813 588 1814 592
rect 2170 588 2171 592
rect 3958 588 3966 591
rect 374 568 410 571
rect 1386 568 1387 572
rect 1794 568 1801 571
rect 3130 568 3131 572
rect 3970 568 4001 571
rect 4326 568 4353 571
rect 598 558 617 561
rect 1158 548 1161 558
rect 1398 558 1414 561
rect 2226 558 2230 562
rect 1514 548 1521 551
rect 1550 548 1558 551
rect 1642 548 1649 551
rect 1850 548 1857 551
rect 1870 548 1878 551
rect 1906 548 1913 551
rect 2090 548 2097 551
rect 2126 548 2145 551
rect 2162 548 2169 551
rect 2270 551 2273 561
rect 2394 558 2398 562
rect 3142 558 3153 561
rect 3550 558 3561 561
rect 2270 548 2289 551
rect 2318 548 2326 551
rect 3070 548 3081 551
rect 3302 548 3310 551
rect 78 538 81 548
rect 174 541 177 548
rect 166 538 177 541
rect 1110 538 1118 541
rect 1694 538 1705 541
rect 1734 538 1753 541
rect 1862 538 1881 541
rect 2294 541 2297 548
rect 2294 538 2313 541
rect 2806 538 2833 541
rect 3102 538 3110 541
rect 3274 538 3289 541
rect 3522 538 3529 541
rect 3606 538 3614 541
rect 3850 538 3857 541
rect 1878 532 1881 538
rect 2054 532 2058 534
rect 1090 528 1102 531
rect 1838 528 1846 531
rect 2198 528 2206 531
rect 3270 528 3273 538
rect 2034 518 2035 522
rect 2698 518 2699 522
rect 2862 518 2878 521
rect 3322 518 3323 522
rect 3597 518 3598 522
rect 3733 518 3734 522
rect 3789 518 3790 522
rect 3813 518 3814 522
rect 3866 518 3867 522
rect 896 503 898 507
rect 902 503 905 507
rect 909 503 912 507
rect 1928 503 1930 507
rect 1934 503 1937 507
rect 1941 503 1944 507
rect 2952 503 2954 507
rect 2958 503 2961 507
rect 2965 503 2968 507
rect 3976 503 3978 507
rect 3982 503 3985 507
rect 3989 503 3992 507
rect 3554 488 3555 492
rect 4378 488 4385 491
rect 4054 478 4065 481
rect 4150 478 4161 481
rect 4062 472 4065 478
rect 4158 472 4161 478
rect 462 468 470 471
rect 1118 468 1126 471
rect 1678 468 1686 471
rect 2470 468 2478 471
rect 2510 462 2513 471
rect 2778 468 2785 471
rect 2810 468 2817 471
rect 3210 468 3217 471
rect 3294 468 3305 471
rect 3314 468 3329 471
rect 3526 468 3553 471
rect 3742 468 3750 471
rect 3762 468 3769 471
rect 3826 468 3833 471
rect 4310 471 4313 478
rect 4318 471 4322 472
rect 4310 468 4322 471
rect 22 458 41 461
rect 1126 458 1134 461
rect 1478 458 1486 461
rect 1502 458 1510 461
rect 1734 458 1750 461
rect 1794 458 1801 461
rect 1846 458 1865 461
rect 2126 458 2134 461
rect 2370 458 2385 461
rect 2482 458 2497 461
rect 2806 458 2814 461
rect 3074 458 3081 461
rect 3086 458 3094 461
rect 3126 458 3134 461
rect 3274 458 3281 461
rect 3650 458 3657 461
rect 3670 458 3689 461
rect 994 448 998 452
rect 1158 448 1177 451
rect 1422 448 1438 451
rect 1730 448 1734 452
rect 1862 448 1865 458
rect 2354 448 2358 452
rect 2826 448 2830 452
rect 3594 448 3598 452
rect 3606 448 3617 451
rect 3670 448 3673 458
rect 3910 448 3921 451
rect 3974 448 3982 451
rect 4310 442 4313 461
rect 1006 438 1025 441
rect 1146 438 1147 442
rect 2125 438 2126 442
rect 2146 438 2153 441
rect 2170 438 2177 441
rect 4338 438 4353 441
rect 1022 428 1025 438
rect 1778 418 1779 422
rect 3250 418 3251 422
rect 3658 418 3659 422
rect 3802 418 3803 422
rect 3986 418 4001 421
rect 392 403 394 407
rect 398 403 401 407
rect 405 403 408 407
rect 1416 403 1418 407
rect 1422 403 1425 407
rect 1429 403 1432 407
rect 2440 403 2442 407
rect 2446 403 2449 407
rect 2453 403 2456 407
rect 3472 403 3474 407
rect 3478 403 3481 407
rect 3485 403 3488 407
rect 1130 388 1131 392
rect 898 368 899 372
rect 942 371 945 381
rect 910 368 945 371
rect 2517 368 2518 372
rect 3853 368 3854 372
rect 486 358 505 361
rect 930 358 937 361
rect 978 358 982 362
rect 990 358 1009 361
rect 1078 358 1089 361
rect 1242 358 1246 362
rect 1326 358 1345 361
rect 1954 358 1969 361
rect 1974 358 1993 361
rect 2750 358 2758 361
rect 2994 358 2998 362
rect 3290 358 3294 362
rect 22 348 30 351
rect 550 348 569 351
rect 574 348 582 351
rect 586 348 601 351
rect 1102 348 1118 351
rect 1146 348 1153 351
rect 1354 348 1361 351
rect 1582 348 1590 351
rect 2290 348 2297 351
rect 2302 348 2329 351
rect 2406 348 2414 351
rect 2518 348 2545 351
rect 2726 348 2734 351
rect 3306 348 3321 351
rect 3326 348 3334 351
rect 3622 348 3638 351
rect 3734 348 3745 351
rect 3974 348 3982 351
rect 282 338 289 341
rect 582 338 590 341
rect 1230 341 1233 348
rect 1114 338 1121 341
rect 1214 338 1233 341
rect 1374 338 1382 341
rect 1542 338 1558 341
rect 2438 338 2454 341
rect 2726 338 2729 348
rect 3078 338 3086 341
rect 3398 338 3422 341
rect 3674 338 3681 341
rect 3686 338 3697 341
rect 3702 338 3718 341
rect 1886 332 1890 334
rect 1306 328 1308 332
rect 3702 328 3705 338
rect 1498 318 1500 322
rect 896 303 898 307
rect 902 303 905 307
rect 909 303 912 307
rect 1928 303 1930 307
rect 1934 303 1937 307
rect 1941 303 1944 307
rect 2952 303 2954 307
rect 2958 303 2961 307
rect 2965 303 2968 307
rect 3976 303 3978 307
rect 3982 303 3985 307
rect 3989 303 3992 307
rect 1541 288 1542 292
rect 1605 288 1606 292
rect 2293 288 2294 292
rect 1134 278 1145 281
rect 1622 278 1633 281
rect 1134 272 1137 278
rect 1622 272 1625 278
rect 930 268 937 271
rect 1142 268 1161 271
rect 1214 268 1225 271
rect 1498 268 1505 271
rect 1518 268 1526 271
rect 2258 268 2265 271
rect 2358 268 2374 271
rect 2438 268 2446 271
rect 2582 268 2590 271
rect 3334 268 3345 271
rect 3510 268 3537 271
rect 1214 262 1217 268
rect 834 258 849 261
rect 950 258 958 261
rect 1470 261 1473 268
rect 3822 268 3833 271
rect 4290 268 4297 271
rect 1454 258 1473 261
rect 1526 258 1534 261
rect 1590 258 1598 261
rect 2162 258 2177 261
rect 2214 258 2233 261
rect 2238 258 2254 261
rect 2326 258 2345 261
rect 2466 258 2473 261
rect 3050 258 3057 261
rect 3358 258 3366 261
rect 3398 258 3406 261
rect 3430 258 3438 261
rect 3654 258 3662 261
rect 3694 258 3702 261
rect 3906 258 3913 261
rect 4030 258 4038 261
rect 1210 248 1217 251
rect 1326 248 1345 251
rect 2054 248 2073 251
rect 2078 248 2086 251
rect 2190 248 2209 251
rect 2214 248 2217 258
rect 2326 248 2329 258
rect 2426 248 2430 252
rect 2513 248 2518 252
rect 2558 248 2569 251
rect 3714 248 3718 252
rect 1190 242 1194 244
rect 866 238 867 242
rect 1254 242 1258 244
rect 1310 238 1318 241
rect 1406 238 1446 241
rect 2149 238 2150 242
rect 3978 238 3985 241
rect 894 228 897 238
rect 2042 228 2043 232
rect 373 218 374 222
rect 2178 218 2179 222
rect 2546 218 2547 222
rect 3653 218 3654 222
rect 3749 218 3750 222
rect 392 203 394 207
rect 398 203 401 207
rect 405 203 408 207
rect 1416 203 1418 207
rect 1422 203 1425 207
rect 1429 203 1432 207
rect 2440 203 2442 207
rect 2446 203 2449 207
rect 2453 203 2456 207
rect 3472 203 3474 207
rect 3478 203 3481 207
rect 3485 203 3488 207
rect 1122 188 1123 192
rect 4285 188 4286 192
rect 834 168 835 172
rect 1010 168 1011 172
rect 1150 171 1153 181
rect 1330 178 1331 182
rect 2613 178 2614 182
rect 1134 168 1153 171
rect 1234 168 1241 171
rect 1266 168 1267 172
rect 1486 168 1494 171
rect 2130 168 2131 172
rect 978 158 982 162
rect 1042 158 1046 162
rect 366 148 401 151
rect 582 148 601 151
rect 782 148 801 151
rect 858 148 865 151
rect 1182 148 1198 151
rect 1290 148 1297 151
rect 1322 148 1329 151
rect 1502 151 1506 154
rect 1502 148 1521 151
rect 1854 151 1858 152
rect 1854 148 1873 151
rect 1894 148 1910 151
rect 2058 148 2065 151
rect 2166 151 2169 161
rect 2590 158 2601 161
rect 2166 148 2185 151
rect 2526 148 2534 151
rect 2758 151 2761 161
rect 2742 148 2761 151
rect 3614 148 3617 158
rect 3914 158 3918 162
rect 4006 148 4014 151
rect 1386 138 1396 141
rect 1534 141 1537 148
rect 1534 138 1545 141
rect 1830 141 1833 148
rect 1822 138 1833 141
rect 1894 141 1897 148
rect 1886 138 1897 141
rect 1934 138 1950 141
rect 1982 138 1993 141
rect 2086 138 2089 148
rect 2230 141 2233 148
rect 2222 138 2233 141
rect 2246 138 2265 141
rect 2438 138 2454 141
rect 2486 138 2513 141
rect 2518 138 2537 141
rect 2658 138 2673 141
rect 2686 138 2705 141
rect 3054 141 3057 148
rect 3046 138 3057 141
rect 3422 138 3430 141
rect 3970 138 3993 141
rect 4014 138 4033 141
rect 4294 138 4302 141
rect 1370 128 1374 132
rect 2670 128 2673 138
rect 3866 128 3873 131
rect 1482 118 1484 122
rect 2162 118 2163 122
rect 2642 118 2643 122
rect 896 103 898 107
rect 902 103 905 107
rect 909 103 912 107
rect 1928 103 1930 107
rect 1934 103 1937 107
rect 1941 103 1944 107
rect 2952 103 2954 107
rect 2958 103 2961 107
rect 2965 103 2968 107
rect 3976 103 3978 107
rect 3982 103 3985 107
rect 3989 103 3992 107
rect 1338 88 1339 92
rect 1410 88 1411 92
rect 2045 88 2046 92
rect 2141 88 2142 92
rect 2317 88 2318 92
rect 2405 88 2406 92
rect 4332 88 4334 92
rect 1114 78 1118 82
rect 2442 78 2449 81
rect 1086 68 1097 71
rect 2014 68 2025 71
rect 2230 68 2238 71
rect 2702 68 2721 71
rect 2726 68 2753 71
rect 2766 68 2774 71
rect 2990 71 2993 78
rect 2982 68 2993 71
rect 3606 71 3609 78
rect 3542 68 3553 71
rect 3574 68 3593 71
rect 3606 68 3625 71
rect 3970 68 3985 71
rect 1086 62 1089 68
rect 46 58 65 61
rect 642 58 649 61
rect 934 58 953 61
rect 1046 58 1065 61
rect 1662 58 1665 68
rect 2014 62 2017 68
rect 1970 58 1993 61
rect 1998 58 2006 61
rect 2210 58 2214 61
rect 2362 58 2369 61
rect 2638 58 2646 61
rect 3038 58 3041 68
rect 3550 62 3553 68
rect 3182 58 3190 61
rect 626 48 630 52
rect 858 48 862 52
rect 2658 48 2662 52
rect 3666 48 3670 52
rect 1086 42 1090 44
rect 1342 42 1346 44
rect 1390 41 1394 44
rect 1390 38 1398 41
rect 1414 41 1418 44
rect 1414 38 1430 41
rect 2142 38 2150 41
rect 390 18 406 21
rect 392 3 394 7
rect 398 3 401 7
rect 405 3 408 7
rect 1416 3 1418 7
rect 1422 3 1425 7
rect 1429 3 1432 7
rect 2440 3 2442 7
rect 2446 3 2449 7
rect 2453 3 2456 7
rect 3472 3 3474 7
rect 3478 3 3481 7
rect 3485 3 3488 7
<< m2contact >>
rect 898 3103 902 3107
rect 905 3103 909 3107
rect 1930 3103 1934 3107
rect 1937 3103 1941 3107
rect 2954 3103 2958 3107
rect 2961 3103 2965 3107
rect 3978 3103 3982 3107
rect 3985 3103 3989 3107
rect 646 3088 650 3092
rect 694 3088 698 3092
rect 1734 3088 1738 3092
rect 1758 3088 1762 3092
rect 1766 3088 1770 3092
rect 1806 3088 1810 3092
rect 2022 3088 2026 3092
rect 2046 3088 2050 3092
rect 3854 3088 3858 3092
rect 230 3078 234 3082
rect 454 3078 458 3082
rect 614 3078 618 3082
rect 6 3068 10 3072
rect 70 3068 74 3072
rect 78 3068 82 3072
rect 214 3068 218 3072
rect 438 3068 442 3072
rect 550 3068 554 3072
rect 566 3068 570 3072
rect 606 3068 610 3072
rect 638 3078 642 3082
rect 654 3078 658 3082
rect 814 3078 818 3082
rect 950 3078 954 3082
rect 1038 3078 1042 3082
rect 1358 3078 1362 3082
rect 1622 3078 1626 3082
rect 1894 3078 1898 3082
rect 2174 3078 2178 3082
rect 2510 3078 2514 3082
rect 2830 3078 2834 3082
rect 3014 3078 3018 3082
rect 3190 3078 3194 3082
rect 3366 3078 3370 3082
rect 3550 3078 3554 3082
rect 3670 3078 3674 3082
rect 3718 3078 3722 3082
rect 3846 3078 3850 3082
rect 4094 3078 4098 3082
rect 4262 3078 4266 3082
rect 4294 3078 4298 3082
rect 678 3068 682 3072
rect 702 3068 706 3072
rect 718 3068 722 3072
rect 734 3068 738 3072
rect 782 3068 786 3072
rect 798 3068 802 3072
rect 838 3068 842 3072
rect 1054 3068 1058 3072
rect 1198 3068 1202 3072
rect 1270 3068 1274 3072
rect 1342 3068 1346 3072
rect 1534 3068 1538 3072
rect 1606 3068 1610 3072
rect 1878 3068 1882 3072
rect 2086 3068 2090 3072
rect 2190 3068 2194 3072
rect 2326 3068 2330 3072
rect 2334 3068 2338 3072
rect 2398 3068 2402 3072
rect 2526 3068 2530 3072
rect 2662 3068 2666 3072
rect 2670 3068 2674 3072
rect 2846 3068 2850 3072
rect 2998 3068 3002 3072
rect 3174 3068 3178 3072
rect 3350 3068 3354 3072
rect 3518 3068 3522 3072
rect 3614 3068 3618 3072
rect 3646 3068 3650 3072
rect 3654 3068 3658 3072
rect 3670 3068 3674 3072
rect 3686 3068 3690 3072
rect 3702 3068 3706 3072
rect 3750 3068 3754 3072
rect 3766 3068 3770 3072
rect 270 3058 274 3062
rect 311 3058 315 3062
rect 350 3058 354 3062
rect 494 3058 498 3062
rect 558 3058 562 3062
rect 598 3058 602 3062
rect 614 3058 618 3062
rect 654 3058 658 3062
rect 670 3058 674 3062
rect 710 3058 714 3062
rect 830 3058 834 3062
rect 846 3058 850 3062
rect 878 3058 882 3062
rect 926 3058 930 3062
rect 998 3058 1002 3062
rect 1150 3058 1154 3062
rect 1294 3058 1298 3062
rect 1398 3058 1402 3062
rect 1662 3058 1666 3062
rect 1742 3058 1746 3062
rect 1782 3058 1786 3062
rect 1790 3058 1794 3062
rect 1838 3058 1842 3062
rect 2030 3058 2034 3062
rect 2054 3058 2058 3062
rect 2134 3058 2138 3062
rect 2470 3058 2474 3062
rect 2894 3058 2898 3062
rect 2958 3058 2962 3062
rect 3126 3058 3130 3062
rect 3134 3058 3138 3062
rect 3230 3058 3234 3062
rect 3302 3058 3306 3062
rect 3494 3058 3498 3062
rect 3526 3058 3530 3062
rect 3550 3058 3554 3062
rect 3574 3058 3578 3062
rect 3614 3058 3618 3062
rect 3694 3058 3698 3062
rect 3742 3058 3746 3062
rect 3766 3058 3770 3062
rect 3790 3058 3794 3062
rect 3862 3068 3866 3072
rect 3910 3068 3914 3072
rect 3958 3068 3962 3072
rect 3966 3068 3970 3072
rect 4078 3068 4082 3072
rect 4102 3068 4106 3072
rect 4142 3068 4146 3072
rect 4206 3068 4210 3072
rect 4230 3068 4234 3072
rect 4246 3068 4250 3072
rect 4278 3068 4282 3072
rect 3822 3058 3826 3062
rect 3870 3058 3874 3062
rect 3886 3058 3890 3062
rect 158 3048 162 3052
rect 182 3050 186 3054
rect 334 3048 338 3052
rect 390 3048 394 3052
rect 582 3048 586 3052
rect 694 3048 698 3052
rect 726 3048 730 3052
rect 750 3048 754 3052
rect 790 3048 794 3052
rect 862 3048 866 3052
rect 942 3048 946 3052
rect 950 3048 954 3052
rect 1102 3048 1106 3052
rect 1134 3048 1138 3052
rect 1294 3048 1298 3052
rect 1558 3048 1562 3052
rect 1830 3048 1834 3052
rect 2222 3050 2226 3054
rect 2558 3050 2562 3054
rect 2606 3048 2610 3052
rect 2878 3050 2882 3054
rect 2966 3050 2970 3054
rect 3142 3050 3146 3054
rect 3302 3048 3306 3052
rect 3502 3048 3506 3052
rect 3582 3048 3586 3052
rect 3590 3048 3594 3052
rect 3622 3048 3626 3052
rect 3670 3048 3674 3052
rect 3758 3048 3762 3052
rect 3774 3048 3778 3052
rect 3790 3048 3794 3052
rect 3814 3048 3818 3052
rect 1262 3038 1266 3042
rect 3502 3038 3506 3042
rect 3518 3038 3522 3042
rect 3566 3038 3570 3042
rect 3830 3038 3834 3042
rect 3886 3038 3890 3042
rect 3926 3058 3930 3062
rect 3950 3058 3954 3062
rect 3990 3058 3994 3062
rect 4014 3058 4018 3062
rect 4038 3058 4042 3062
rect 4054 3058 4058 3062
rect 4118 3058 4122 3062
rect 4150 3058 4154 3062
rect 4182 3058 4186 3062
rect 4230 3058 4234 3062
rect 4238 3058 4242 3062
rect 4270 3058 4274 3062
rect 4310 3058 4314 3062
rect 4390 3058 4394 3062
rect 3902 3048 3906 3052
rect 3926 3048 3930 3052
rect 3990 3048 3994 3052
rect 4030 3048 4034 3052
rect 4110 3048 4114 3052
rect 4166 3048 4170 3052
rect 4174 3048 4178 3052
rect 4206 3048 4210 3052
rect 4302 3048 4306 3052
rect 3998 3038 4002 3042
rect 4022 3038 4026 3042
rect 4126 3038 4130 3042
rect 4190 3038 4194 3042
rect 4318 3038 4322 3042
rect 270 3027 274 3031
rect 494 3027 498 3031
rect 534 3028 538 3032
rect 998 3027 1002 3031
rect 2222 3027 2226 3031
rect 2966 3027 2970 3031
rect 3094 3028 3098 3032
rect 3606 3028 3610 3032
rect 134 3018 138 3022
rect 822 3018 826 3022
rect 1182 3018 1186 3022
rect 1206 3018 1210 3022
rect 1294 3018 1298 3022
rect 1438 3018 1442 3022
rect 1478 3018 1482 3022
rect 1558 3018 1562 3022
rect 1830 3018 1834 3022
rect 2094 3018 2098 3022
rect 2270 3018 2274 3022
rect 2342 3018 2346 3022
rect 2430 3018 2434 3022
rect 2558 3018 2562 3022
rect 2726 3018 2730 3022
rect 2750 3018 2754 3022
rect 2878 3018 2882 3022
rect 3142 3018 3146 3022
rect 3270 3018 3274 3022
rect 3302 3018 3306 3022
rect 3446 3018 3450 3022
rect 3494 3018 3498 3022
rect 3574 3018 3578 3022
rect 3638 3018 3642 3022
rect 3742 3018 3746 3022
rect 3822 3018 3826 3022
rect 3878 3018 3882 3022
rect 4046 3018 4050 3022
rect 4118 3018 4122 3022
rect 4150 3018 4154 3022
rect 4198 3018 4202 3022
rect 4262 3018 4266 3022
rect 4294 3018 4298 3022
rect 4326 3018 4330 3022
rect 4342 3018 4346 3022
rect 394 3003 398 3007
rect 401 3003 405 3007
rect 1418 3003 1422 3007
rect 1425 3003 1429 3007
rect 2442 3003 2446 3007
rect 2449 3003 2453 3007
rect 3474 3003 3478 3007
rect 3481 3003 3485 3007
rect 1230 2988 1234 2992
rect 1630 2988 1634 2992
rect 1798 2988 1802 2992
rect 1942 2988 1946 2992
rect 2070 2988 2074 2992
rect 2086 2988 2090 2992
rect 2230 2988 2234 2992
rect 2606 2988 2610 2992
rect 2854 2988 2858 2992
rect 3054 2988 3058 2992
rect 3086 2988 3090 2992
rect 3166 2988 3170 2992
rect 3198 2988 3202 2992
rect 3758 2988 3762 2992
rect 3766 2988 3770 2992
rect 3998 2988 4002 2992
rect 4166 2988 4170 2992
rect 4246 2988 4250 2992
rect 4294 2988 4298 2992
rect 4366 2988 4370 2992
rect 110 2978 114 2982
rect 246 2978 250 2982
rect 782 2978 786 2982
rect 1142 2978 1146 2982
rect 1534 2978 1538 2982
rect 3246 2979 3250 2983
rect 3438 2978 3442 2982
rect 2574 2968 2578 2972
rect 2806 2968 2810 2972
rect 2902 2968 2906 2972
rect 3446 2968 3450 2972
rect 3566 2968 3570 2972
rect 3718 2968 3722 2972
rect 3750 2968 3754 2972
rect 3806 2968 3810 2972
rect 4110 2968 4114 2972
rect 4118 2968 4122 2972
rect 4142 2968 4146 2972
rect 4174 2968 4178 2972
rect 4374 2968 4378 2972
rect 158 2958 162 2962
rect 214 2956 218 2960
rect 622 2958 626 2962
rect 830 2958 834 2962
rect 862 2958 866 2962
rect 950 2958 954 2962
rect 974 2958 978 2962
rect 998 2958 1002 2962
rect 1174 2956 1178 2960
rect 1230 2958 1234 2962
rect 1510 2958 1514 2962
rect 110 2948 114 2952
rect 246 2948 250 2952
rect 343 2948 347 2952
rect 438 2948 442 2952
rect 478 2948 482 2952
rect 542 2948 546 2952
rect 590 2948 594 2952
rect 622 2948 626 2952
rect 670 2948 674 2952
rect 685 2948 689 2952
rect 782 2948 786 2952
rect 870 2948 874 2952
rect 878 2948 882 2952
rect 998 2948 1002 2952
rect 1030 2948 1034 2952
rect 1142 2948 1146 2952
rect 1238 2948 1242 2952
rect 1398 2948 1402 2952
rect 1414 2948 1418 2952
rect 1454 2948 1458 2952
rect 1462 2948 1466 2952
rect 1470 2948 1474 2952
rect 1494 2948 1498 2952
rect 1582 2958 1586 2962
rect 1630 2958 1634 2962
rect 1942 2958 1946 2962
rect 2230 2958 2234 2962
rect 2270 2958 2274 2962
rect 1534 2948 1538 2952
rect 1638 2948 1642 2952
rect 1838 2948 1842 2952
rect 2054 2948 2058 2952
rect 2126 2948 2130 2952
rect 2214 2948 2218 2952
rect 2606 2958 2610 2962
rect 2758 2958 2762 2962
rect 2822 2958 2826 2962
rect 2870 2958 2874 2962
rect 3142 2958 3146 2962
rect 2294 2948 2298 2952
rect 2326 2948 2330 2952
rect 2566 2948 2570 2952
rect 2606 2948 2610 2952
rect 110 2938 114 2942
rect 246 2938 250 2942
rect 358 2938 362 2942
rect 374 2938 378 2942
rect 558 2938 562 2942
rect 606 2938 610 2942
rect 622 2938 626 2942
rect 654 2938 658 2942
rect 782 2938 786 2942
rect 886 2938 890 2942
rect 926 2938 930 2942
rect 942 2938 946 2942
rect 958 2938 962 2942
rect 974 2938 978 2942
rect 1006 2938 1010 2942
rect 1142 2938 1146 2942
rect 1278 2938 1282 2942
rect 1390 2938 1394 2942
rect 1406 2938 1410 2942
rect 1422 2938 1426 2942
rect 1478 2938 1482 2942
rect 1486 2938 1490 2942
rect 1542 2938 1546 2942
rect 1558 2938 1562 2942
rect 1598 2938 1602 2942
rect 1678 2938 1682 2942
rect 1894 2938 1898 2942
rect 1966 2938 1970 2942
rect 2182 2938 2186 2942
rect 2254 2938 2258 2942
rect 2302 2938 2306 2942
rect 2398 2938 2402 2942
rect 2470 2938 2474 2942
rect 2558 2938 2562 2942
rect 2654 2938 2658 2942
rect 2782 2938 2786 2942
rect 2798 2948 2802 2952
rect 2878 2948 2882 2952
rect 2974 2948 2978 2952
rect 3070 2948 3074 2952
rect 3102 2948 3106 2952
rect 3182 2958 3186 2962
rect 3246 2956 3250 2960
rect 3430 2958 3434 2962
rect 3486 2958 3490 2962
rect 3582 2958 3586 2962
rect 3702 2958 3706 2962
rect 3734 2958 3738 2962
rect 3902 2958 3906 2962
rect 3942 2958 3946 2962
rect 3982 2958 3986 2962
rect 4038 2958 4042 2962
rect 4102 2958 4106 2962
rect 4158 2958 4162 2962
rect 4190 2958 4194 2962
rect 4214 2958 4218 2962
rect 4222 2958 4226 2962
rect 4262 2958 4266 2962
rect 4350 2958 4354 2962
rect 4358 2958 4362 2962
rect 3166 2948 3170 2952
rect 3198 2948 3202 2952
rect 3230 2948 3234 2952
rect 3334 2948 3338 2952
rect 3422 2948 3426 2952
rect 3438 2948 3442 2952
rect 3478 2948 3482 2952
rect 3566 2948 3570 2952
rect 3590 2948 3594 2952
rect 3614 2948 3618 2952
rect 3662 2948 3666 2952
rect 3670 2948 3674 2952
rect 3710 2948 3714 2952
rect 3742 2948 3746 2952
rect 3790 2948 3794 2952
rect 3846 2948 3850 2952
rect 3886 2948 3890 2952
rect 3998 2948 4002 2952
rect 4014 2948 4018 2952
rect 4030 2948 4034 2952
rect 4062 2948 4066 2952
rect 4094 2948 4098 2952
rect 4110 2948 4114 2952
rect 4150 2948 4154 2952
rect 4182 2948 4186 2952
rect 4262 2948 4266 2952
rect 4278 2948 4282 2952
rect 4326 2948 4330 2952
rect 4350 2948 4354 2952
rect 4366 2948 4370 2952
rect 2838 2938 2842 2942
rect 2846 2938 2850 2942
rect 2886 2938 2890 2942
rect 2910 2938 2914 2942
rect 2998 2938 3002 2942
rect 3126 2938 3130 2942
rect 3174 2938 3178 2942
rect 3206 2938 3210 2942
rect 3278 2938 3282 2942
rect 3406 2938 3410 2942
rect 3502 2938 3506 2942
rect 3550 2938 3554 2942
rect 3558 2938 3562 2942
rect 3622 2938 3626 2942
rect 3678 2938 3682 2942
rect 3854 2938 3858 2942
rect 3926 2938 3930 2942
rect 3958 2938 3962 2942
rect 4006 2938 4010 2942
rect 4054 2938 4058 2942
rect 4086 2938 4090 2942
rect 4150 2938 4154 2942
rect 4198 2938 4202 2942
rect 4238 2938 4242 2942
rect 4286 2938 4290 2942
rect 4310 2938 4314 2942
rect 6 2928 10 2932
rect 94 2928 98 2932
rect 262 2928 266 2932
rect 382 2928 386 2932
rect 414 2928 418 2932
rect 422 2928 426 2932
rect 446 2928 450 2932
rect 566 2928 570 2932
rect 630 2928 634 2932
rect 654 2928 658 2932
rect 766 2928 770 2932
rect 854 2928 858 2932
rect 902 2928 906 2932
rect 1038 2928 1042 2932
rect 1126 2928 1130 2932
rect 1294 2928 1298 2932
rect 1550 2928 1554 2932
rect 1574 2928 1578 2932
rect 1606 2928 1610 2932
rect 1694 2928 1698 2932
rect 1878 2928 1882 2932
rect 2166 2928 2170 2932
rect 2582 2928 2586 2932
rect 2670 2928 2674 2932
rect 2766 2928 2770 2932
rect 2814 2928 2818 2932
rect 2902 2928 2906 2932
rect 3118 2928 3122 2932
rect 3294 2928 3298 2932
rect 3390 2928 3394 2932
rect 3406 2928 3410 2932
rect 3422 2928 3426 2932
rect 3494 2928 3498 2932
rect 3638 2928 3642 2932
rect 3694 2928 3698 2932
rect 3766 2928 3770 2932
rect 3814 2928 3818 2932
rect 3846 2928 3850 2932
rect 3854 2928 3858 2932
rect 4030 2928 4034 2932
rect 4038 2928 4042 2932
rect 4070 2928 4074 2932
rect 4078 2928 4082 2932
rect 4254 2928 4258 2932
rect 4318 2928 4322 2932
rect 430 2918 434 2922
rect 470 2918 474 2922
rect 494 2918 498 2922
rect 550 2918 554 2922
rect 566 2918 570 2922
rect 662 2918 666 2922
rect 974 2918 978 2922
rect 1374 2918 1378 2922
rect 1774 2918 1778 2922
rect 2038 2918 2042 2922
rect 2278 2918 2282 2922
rect 2342 2918 2346 2922
rect 2414 2918 2418 2922
rect 2750 2918 2754 2922
rect 3054 2918 3058 2922
rect 3110 2918 3114 2922
rect 3374 2918 3378 2922
rect 3534 2918 3538 2922
rect 3630 2918 3634 2922
rect 3686 2918 3690 2922
rect 3718 2918 3722 2922
rect 3918 2918 3922 2922
rect 4206 2918 4210 2922
rect 4230 2918 4234 2922
rect 898 2903 902 2907
rect 905 2903 909 2907
rect 1930 2903 1934 2907
rect 1937 2903 1941 2907
rect 2954 2903 2958 2907
rect 2961 2903 2965 2907
rect 3978 2903 3982 2907
rect 3985 2903 3989 2907
rect 838 2888 842 2892
rect 870 2888 874 2892
rect 926 2888 930 2892
rect 982 2888 986 2892
rect 1006 2888 1010 2892
rect 1046 2888 1050 2892
rect 1406 2888 1410 2892
rect 1430 2888 1434 2892
rect 1566 2888 1570 2892
rect 1582 2888 1586 2892
rect 2030 2888 2034 2892
rect 2086 2888 2090 2892
rect 2630 2888 2634 2892
rect 2942 2888 2946 2892
rect 3182 2888 3186 2892
rect 3206 2888 3210 2892
rect 3502 2888 3506 2892
rect 3558 2888 3562 2892
rect 3582 2888 3586 2892
rect 3702 2888 3706 2892
rect 3782 2888 3786 2892
rect 3854 2888 3858 2892
rect 4134 2888 4138 2892
rect 4166 2888 4170 2892
rect 4238 2888 4242 2892
rect 22 2878 26 2882
rect 174 2878 178 2882
rect 270 2878 274 2882
rect 358 2878 362 2882
rect 558 2878 562 2882
rect 566 2878 570 2882
rect 606 2878 610 2882
rect 630 2878 634 2882
rect 750 2878 754 2882
rect 918 2878 922 2882
rect 1270 2878 1274 2882
rect 1406 2878 1410 2882
rect 1422 2878 1426 2882
rect 30 2868 34 2872
rect 102 2868 106 2872
rect 190 2868 194 2872
rect 238 2868 242 2872
rect 254 2868 258 2872
rect 342 2868 346 2872
rect 470 2868 474 2872
rect 502 2868 506 2872
rect 518 2868 522 2872
rect 646 2868 650 2872
rect 654 2868 658 2872
rect 766 2868 770 2872
rect 854 2868 858 2872
rect 950 2868 954 2872
rect 958 2868 962 2872
rect 990 2868 994 2872
rect 1038 2868 1042 2872
rect 1070 2868 1074 2872
rect 1078 2868 1082 2872
rect 1182 2868 1186 2872
rect 1254 2868 1258 2872
rect 1382 2868 1386 2872
rect 1438 2868 1442 2872
rect 1542 2868 1546 2872
rect 1638 2868 1642 2872
rect 1742 2868 1746 2872
rect 1950 2878 1954 2882
rect 2046 2878 2050 2882
rect 2174 2878 2178 2882
rect 2310 2878 2314 2882
rect 2422 2878 2426 2882
rect 2566 2878 2570 2882
rect 2750 2878 2754 2882
rect 2838 2878 2842 2882
rect 2934 2878 2938 2882
rect 2982 2878 2986 2882
rect 3078 2878 3082 2882
rect 3366 2878 3370 2882
rect 3518 2878 3522 2882
rect 3550 2878 3554 2882
rect 3630 2878 3634 2882
rect 3766 2878 3770 2882
rect 3862 2878 3866 2882
rect 3886 2878 3890 2882
rect 3910 2878 3914 2882
rect 3990 2878 3994 2882
rect 4030 2878 4034 2882
rect 4094 2878 4098 2882
rect 4126 2878 4130 2882
rect 4238 2878 4242 2882
rect 1934 2868 1938 2872
rect 2158 2868 2162 2872
rect 2318 2868 2322 2872
rect 2334 2868 2338 2872
rect 2438 2868 2442 2872
rect 2526 2868 2530 2872
rect 2542 2868 2546 2872
rect 2582 2868 2586 2872
rect 2614 2868 2618 2872
rect 2662 2868 2666 2872
rect 2766 2868 2770 2872
rect 2846 2868 2850 2872
rect 2862 2868 2866 2872
rect 2950 2868 2954 2872
rect 3094 2868 3098 2872
rect 3166 2868 3170 2872
rect 3198 2868 3202 2872
rect 3214 2868 3218 2872
rect 3270 2868 3274 2872
rect 3278 2868 3282 2872
rect 3350 2868 3354 2872
rect 3462 2868 3466 2872
rect 3510 2868 3514 2872
rect 3550 2868 3554 2872
rect 3574 2868 3578 2872
rect 3598 2868 3602 2872
rect 6 2858 10 2862
rect 230 2858 234 2862
rect 246 2858 250 2862
rect 270 2858 274 2862
rect 398 2858 402 2862
rect 478 2858 482 2862
rect 542 2858 546 2862
rect 590 2858 594 2862
rect 622 2858 626 2862
rect 662 2858 666 2862
rect 710 2858 714 2862
rect 870 2858 874 2862
rect 902 2858 906 2862
rect 942 2858 946 2862
rect 966 2858 970 2862
rect 1062 2858 1066 2862
rect 1206 2858 1210 2862
rect 1366 2858 1370 2862
rect 1446 2858 1450 2862
rect 1470 2858 1474 2862
rect 1542 2858 1546 2862
rect 1654 2858 1658 2862
rect 1750 2858 1754 2862
rect 1782 2858 1786 2862
rect 1790 2858 1794 2862
rect 1814 2858 1818 2862
rect 1846 2858 1850 2862
rect 1886 2858 1890 2862
rect 2070 2858 2074 2862
rect 2102 2858 2106 2862
rect 2214 2858 2218 2862
rect 2262 2858 2266 2862
rect 2286 2858 2290 2862
rect 2382 2858 2386 2862
rect 2478 2858 2482 2862
rect 2534 2858 2538 2862
rect 2550 2858 2554 2862
rect 2590 2858 2594 2862
rect 2606 2858 2610 2862
rect 2654 2858 2658 2862
rect 2814 2858 2818 2862
rect 2854 2858 2858 2862
rect 3134 2858 3138 2862
rect 3190 2858 3194 2862
rect 3222 2858 3226 2862
rect 3238 2858 3242 2862
rect 3254 2858 3258 2862
rect 3262 2858 3266 2862
rect 3318 2858 3322 2862
rect 3486 2858 3490 2862
rect 3502 2858 3506 2862
rect 3542 2858 3546 2862
rect 3566 2858 3570 2862
rect 3598 2858 3602 2862
rect 3622 2858 3626 2862
rect 3646 2858 3650 2862
rect 3662 2858 3666 2862
rect 3678 2858 3682 2862
rect 3694 2868 3698 2872
rect 3710 2868 3714 2872
rect 3806 2868 3810 2872
rect 3854 2868 3858 2872
rect 3926 2868 3930 2872
rect 3966 2868 3970 2872
rect 4006 2868 4010 2872
rect 4014 2868 4018 2872
rect 4070 2868 4074 2872
rect 4126 2868 4130 2872
rect 4142 2868 4146 2872
rect 4198 2868 4202 2872
rect 4206 2868 4210 2872
rect 4238 2868 4242 2872
rect 4270 2868 4274 2872
rect 4318 2868 4322 2872
rect 4334 2868 4338 2872
rect 3766 2858 3770 2862
rect 3798 2858 3802 2862
rect 3846 2858 3850 2862
rect 3886 2858 3890 2862
rect 3934 2858 3938 2862
rect 3942 2858 3946 2862
rect 3958 2858 3962 2862
rect 4046 2858 4050 2862
rect 4110 2858 4114 2862
rect 4142 2858 4146 2862
rect 4246 2858 4250 2862
rect 4294 2858 4298 2862
rect 4318 2858 4322 2862
rect 4350 2858 4354 2862
rect 4382 2858 4386 2862
rect 214 2848 218 2852
rect 310 2850 314 2854
rect 494 2848 498 2852
rect 502 2848 506 2852
rect 574 2848 578 2852
rect 630 2848 634 2852
rect 814 2848 818 2852
rect 838 2848 842 2852
rect 870 2848 874 2852
rect 926 2848 930 2852
rect 982 2848 986 2852
rect 1046 2848 1050 2852
rect 1222 2850 1226 2854
rect 1406 2848 1410 2852
rect 1670 2848 1674 2852
rect 1766 2848 1770 2852
rect 1902 2850 1906 2854
rect 2086 2848 2090 2852
rect 2126 2850 2130 2854
rect 2270 2848 2274 2852
rect 2470 2850 2474 2854
rect 2622 2848 2626 2852
rect 2630 2848 2634 2852
rect 2814 2848 2818 2852
rect 3126 2850 3130 2854
rect 3182 2848 3186 2852
rect 3230 2848 3234 2852
rect 3302 2848 3306 2852
rect 3518 2848 3522 2852
rect 3590 2848 3594 2852
rect 3622 2848 3626 2852
rect 3782 2848 3786 2852
rect 3878 2848 3882 2852
rect 3910 2848 3914 2852
rect 3942 2848 3946 2852
rect 3982 2848 3986 2852
rect 4030 2848 4034 2852
rect 4086 2848 4090 2852
rect 4214 2848 4218 2852
rect 4310 2848 4314 2852
rect 4366 2848 4370 2852
rect 534 2838 538 2842
rect 854 2838 858 2842
rect 1662 2838 1666 2842
rect 3662 2838 3666 2842
rect 3894 2838 3898 2842
rect 4038 2838 4042 2842
rect 398 2827 402 2831
rect 710 2827 714 2831
rect 1222 2827 1226 2831
rect 1374 2828 1378 2832
rect 1854 2828 1858 2832
rect 1902 2827 1906 2831
rect 2470 2827 2474 2831
rect 3126 2827 3130 2831
rect 4046 2828 4050 2832
rect 14 2818 18 2822
rect 86 2818 90 2822
rect 158 2818 162 2822
rect 438 2818 442 2822
rect 478 2818 482 2822
rect 526 2818 530 2822
rect 590 2818 594 2822
rect 1126 2818 1130 2822
rect 1486 2818 1490 2822
rect 1646 2818 1650 2822
rect 1686 2818 1690 2822
rect 2126 2818 2130 2822
rect 2254 2818 2258 2822
rect 2342 2818 2346 2822
rect 2670 2818 2674 2822
rect 2814 2818 2818 2822
rect 2918 2818 2922 2822
rect 2998 2818 3002 2822
rect 3302 2818 3306 2822
rect 3446 2818 3450 2822
rect 3742 2818 3746 2822
rect 394 2803 398 2807
rect 401 2803 405 2807
rect 1418 2803 1422 2807
rect 1425 2803 1429 2807
rect 2442 2803 2446 2807
rect 2449 2803 2453 2807
rect 3474 2803 3478 2807
rect 3481 2803 3485 2807
rect 62 2788 66 2792
rect 198 2788 202 2792
rect 558 2788 562 2792
rect 582 2788 586 2792
rect 742 2788 746 2792
rect 1214 2788 1218 2792
rect 1246 2788 1250 2792
rect 1462 2788 1466 2792
rect 1518 2788 1522 2792
rect 1662 2788 1666 2792
rect 1702 2788 1706 2792
rect 1718 2788 1722 2792
rect 1862 2788 1866 2792
rect 2054 2788 2058 2792
rect 2086 2788 2090 2792
rect 2462 2788 2466 2792
rect 2494 2788 2498 2792
rect 2606 2788 2610 2792
rect 2654 2788 2658 2792
rect 2766 2788 2770 2792
rect 3446 2788 3450 2792
rect 3502 2788 3506 2792
rect 4206 2788 4210 2792
rect 4286 2788 4290 2792
rect 430 2778 434 2782
rect 686 2778 690 2782
rect 1302 2779 1306 2783
rect 2270 2779 2274 2783
rect 3046 2779 3050 2783
rect 3190 2779 3194 2783
rect 3318 2778 3322 2782
rect 534 2768 538 2772
rect 1446 2768 1450 2772
rect 2094 2768 2098 2772
rect 2558 2768 2562 2772
rect 2630 2768 2634 2772
rect 3094 2768 3098 2772
rect 3438 2768 3442 2772
rect 3454 2768 3458 2772
rect 3798 2768 3802 2772
rect 4198 2768 4202 2772
rect 4318 2768 4322 2772
rect 6 2758 10 2762
rect 22 2758 26 2762
rect 190 2758 194 2762
rect 302 2758 306 2762
rect 486 2758 490 2762
rect 502 2758 506 2762
rect 550 2758 554 2762
rect 598 2758 602 2762
rect 678 2758 682 2762
rect 726 2758 730 2762
rect 30 2748 34 2752
rect 38 2748 42 2752
rect 70 2748 74 2752
rect 102 2748 106 2752
rect 158 2748 162 2752
rect 286 2748 290 2752
rect 318 2748 322 2752
rect 430 2748 434 2752
rect 526 2748 530 2752
rect 574 2748 578 2752
rect 718 2748 722 2752
rect 742 2748 746 2752
rect 758 2748 762 2752
rect 990 2758 994 2762
rect 1214 2758 1218 2762
rect 1302 2756 1306 2760
rect 1662 2758 1666 2762
rect 1670 2758 1674 2762
rect 1862 2758 1866 2762
rect 2054 2758 2058 2762
rect 2078 2758 2082 2762
rect 2206 2758 2210 2762
rect 806 2748 810 2752
rect 822 2748 826 2752
rect 862 2748 866 2752
rect 886 2748 890 2752
rect 910 2748 914 2752
rect 918 2748 922 2752
rect 974 2748 978 2752
rect 1006 2748 1010 2752
rect 1038 2748 1042 2752
rect 1206 2748 1210 2752
rect 1262 2748 1266 2752
rect 1286 2748 1290 2752
rect 1390 2748 1394 2752
rect 1478 2748 1482 2752
rect 1502 2748 1506 2752
rect 1558 2748 1562 2752
rect 2270 2756 2274 2760
rect 2574 2758 2578 2762
rect 2590 2758 2594 2762
rect 2638 2758 2642 2762
rect 2750 2758 2754 2762
rect 2798 2758 2802 2762
rect 2862 2758 2866 2762
rect 3046 2756 3050 2760
rect 3126 2758 3130 2762
rect 3190 2756 3194 2760
rect 3470 2758 3474 2762
rect 3542 2758 3546 2762
rect 3686 2758 3690 2762
rect 3702 2758 3706 2762
rect 3782 2758 3786 2762
rect 3798 2758 3802 2762
rect 3838 2758 3842 2762
rect 3950 2758 3954 2762
rect 4038 2758 4042 2762
rect 1686 2748 1690 2752
rect 1758 2748 1762 2752
rect 1870 2748 1874 2752
rect 2054 2748 2058 2752
rect 2086 2748 2090 2752
rect 2110 2748 2114 2752
rect 2118 2748 2122 2752
rect 2134 2748 2138 2752
rect 2142 2748 2146 2752
rect 2150 2748 2154 2752
rect 2166 2748 2170 2752
rect 2222 2748 2226 2752
rect 2262 2748 2266 2752
rect 2358 2748 2362 2752
rect 2454 2748 2458 2752
rect 2470 2748 2474 2752
rect 2510 2748 2514 2752
rect 2534 2748 2538 2752
rect 2574 2748 2578 2752
rect 2654 2748 2658 2752
rect 2670 2748 2674 2752
rect 2686 2748 2690 2752
rect 2734 2748 2738 2752
rect 2750 2748 2754 2752
rect 2782 2748 2786 2752
rect 2814 2748 2818 2752
rect 2822 2748 2826 2752
rect 2878 2748 2882 2752
rect 2958 2748 2962 2752
rect 3062 2748 3066 2752
rect 3086 2748 3090 2752
rect 3110 2748 3114 2752
rect 3142 2748 3146 2752
rect 3174 2748 3178 2752
rect 3278 2748 3282 2752
rect 3390 2748 3394 2752
rect 3438 2748 3442 2752
rect 3462 2748 3466 2752
rect 3502 2748 3506 2752
rect 3566 2748 3570 2752
rect 3662 2748 3666 2752
rect 3734 2748 3738 2752
rect 3742 2748 3746 2752
rect 3838 2748 3842 2752
rect 3854 2748 3858 2752
rect 3862 2748 3866 2752
rect 3902 2748 3906 2752
rect 3934 2748 3938 2752
rect 3958 2748 3962 2752
rect 3990 2748 3994 2752
rect 4062 2758 4066 2762
rect 4110 2758 4114 2762
rect 4126 2758 4130 2762
rect 4214 2758 4218 2762
rect 4222 2758 4226 2762
rect 4302 2758 4306 2762
rect 4102 2748 4106 2752
rect 4166 2748 4170 2752
rect 4206 2748 4210 2752
rect 4222 2748 4226 2752
rect 4238 2748 4242 2752
rect 30 2738 34 2742
rect 46 2738 50 2742
rect 78 2738 82 2742
rect 94 2738 98 2742
rect 102 2738 106 2742
rect 150 2738 154 2742
rect 174 2738 178 2742
rect 238 2738 242 2742
rect 254 2738 258 2742
rect 278 2738 282 2742
rect 310 2738 314 2742
rect 430 2738 434 2742
rect 502 2738 506 2742
rect 518 2738 522 2742
rect 526 2738 530 2742
rect 574 2738 578 2742
rect 606 2738 610 2742
rect 750 2738 754 2742
rect 782 2738 786 2742
rect 798 2738 802 2742
rect 830 2738 834 2742
rect 854 2738 858 2742
rect 870 2738 874 2742
rect 894 2738 898 2742
rect 982 2738 986 2742
rect 998 2738 1002 2742
rect 1014 2738 1018 2742
rect 1022 2738 1026 2742
rect 1054 2738 1058 2742
rect 1166 2738 1170 2742
rect 1334 2738 1338 2742
rect 1614 2738 1618 2742
rect 1814 2738 1818 2742
rect 2006 2738 2010 2742
rect 2198 2738 2202 2742
rect 2230 2738 2234 2742
rect 2302 2738 2306 2742
rect 2414 2738 2418 2742
rect 2478 2738 2482 2742
rect 2486 2738 2490 2742
rect 2542 2738 2546 2742
rect 2566 2738 2570 2742
rect 2662 2738 2666 2742
rect 2694 2738 2698 2742
rect 2702 2738 2706 2742
rect 2726 2738 2730 2742
rect 2758 2738 2762 2742
rect 2790 2738 2794 2742
rect 2798 2738 2802 2742
rect 2830 2738 2834 2742
rect 2838 2738 2842 2742
rect 2886 2738 2890 2742
rect 3014 2738 3018 2742
rect 3086 2738 3090 2742
rect 3118 2738 3122 2742
rect 3126 2738 3130 2742
rect 3150 2738 3154 2742
rect 3222 2738 3226 2742
rect 3382 2738 3386 2742
rect 3398 2738 3402 2742
rect 3494 2738 3498 2742
rect 3526 2738 3530 2742
rect 3550 2738 3554 2742
rect 3574 2738 3578 2742
rect 3590 2738 3594 2742
rect 3646 2738 3650 2742
rect 3654 2738 3658 2742
rect 3758 2738 3762 2742
rect 3798 2738 3802 2742
rect 3830 2738 3834 2742
rect 3870 2738 3874 2742
rect 3886 2738 3890 2742
rect 3942 2738 3946 2742
rect 4006 2738 4010 2742
rect 4062 2738 4066 2742
rect 4078 2738 4082 2742
rect 4150 2738 4154 2742
rect 4246 2738 4250 2742
rect 4310 2748 4314 2752
rect 4294 2738 4298 2742
rect 4334 2738 4338 2742
rect 4382 2738 4386 2742
rect 62 2728 66 2732
rect 94 2728 98 2732
rect 118 2728 122 2732
rect 166 2728 170 2732
rect 222 2728 226 2732
rect 270 2728 274 2732
rect 414 2728 418 2732
rect 566 2728 570 2732
rect 702 2728 706 2732
rect 774 2728 778 2732
rect 838 2728 842 2732
rect 870 2728 874 2732
rect 902 2728 906 2732
rect 950 2728 954 2732
rect 1022 2728 1026 2732
rect 1150 2728 1154 2732
rect 1350 2728 1354 2732
rect 1598 2728 1602 2732
rect 1798 2728 1802 2732
rect 1990 2728 1994 2732
rect 2318 2728 2322 2732
rect 2526 2728 2530 2732
rect 2558 2728 2562 2732
rect 2598 2728 2602 2732
rect 2622 2728 2626 2732
rect 2686 2728 2690 2732
rect 2718 2728 2722 2732
rect 2750 2728 2754 2732
rect 2998 2728 3002 2732
rect 3238 2728 3242 2732
rect 3406 2728 3410 2732
rect 3422 2728 3426 2732
rect 3590 2728 3594 2732
rect 3710 2728 3714 2732
rect 3774 2728 3778 2732
rect 3830 2728 3834 2732
rect 3870 2728 3874 2732
rect 3982 2728 3986 2732
rect 4126 2728 4130 2732
rect 4254 2728 4258 2732
rect 4270 2728 4274 2732
rect 662 2718 666 2722
rect 846 2718 850 2722
rect 958 2718 962 2722
rect 1046 2718 1050 2722
rect 1430 2718 1434 2722
rect 1910 2718 1914 2722
rect 2398 2718 2402 2722
rect 2430 2718 2434 2722
rect 2710 2718 2714 2722
rect 2846 2718 2850 2722
rect 2918 2718 2922 2722
rect 3366 2718 3370 2722
rect 3582 2718 3586 2722
rect 3630 2718 3634 2722
rect 3702 2718 3706 2722
rect 3718 2718 3722 2722
rect 3750 2718 3754 2722
rect 3918 2718 3922 2722
rect 3974 2718 3978 2722
rect 4054 2718 4058 2722
rect 4086 2718 4090 2722
rect 4134 2718 4138 2722
rect 4182 2718 4186 2722
rect 4318 2718 4322 2722
rect 4350 2718 4354 2722
rect 898 2703 902 2707
rect 905 2703 909 2707
rect 1930 2703 1934 2707
rect 1937 2703 1941 2707
rect 2954 2703 2958 2707
rect 2961 2703 2965 2707
rect 3978 2703 3982 2707
rect 3985 2703 3989 2707
rect 326 2688 330 2692
rect 422 2688 426 2692
rect 534 2688 538 2692
rect 566 2688 570 2692
rect 630 2688 634 2692
rect 806 2688 810 2692
rect 878 2688 882 2692
rect 902 2688 906 2692
rect 1142 2688 1146 2692
rect 1166 2688 1170 2692
rect 1182 2688 1186 2692
rect 1214 2688 1218 2692
rect 1622 2688 1626 2692
rect 1926 2688 1930 2692
rect 2158 2688 2162 2692
rect 2214 2688 2218 2692
rect 2398 2688 2402 2692
rect 2678 2688 2682 2692
rect 2734 2688 2738 2692
rect 2774 2688 2778 2692
rect 3030 2688 3034 2692
rect 3094 2688 3098 2692
rect 3142 2688 3146 2692
rect 3190 2688 3194 2692
rect 3254 2688 3258 2692
rect 3646 2688 3650 2692
rect 3798 2688 3802 2692
rect 4030 2688 4034 2692
rect 4102 2688 4106 2692
rect 86 2678 90 2682
rect 182 2678 186 2682
rect 214 2678 218 2682
rect 390 2678 394 2682
rect 430 2678 434 2682
rect 446 2678 450 2682
rect 726 2678 730 2682
rect 814 2678 818 2682
rect 886 2678 890 2682
rect 950 2678 954 2682
rect 1038 2678 1042 2682
rect 1350 2678 1354 2682
rect 1542 2678 1546 2682
rect 1750 2678 1754 2682
rect 2046 2678 2050 2682
rect 2262 2678 2266 2682
rect 2390 2678 2394 2682
rect 2422 2678 2426 2682
rect 2582 2678 2586 2682
rect 2686 2678 2690 2682
rect 2814 2678 2818 2682
rect 2902 2678 2906 2682
rect 3262 2678 3266 2682
rect 3430 2678 3434 2682
rect 3582 2678 3586 2682
rect 3614 2678 3618 2682
rect 70 2668 74 2672
rect 214 2668 218 2672
rect 230 2668 234 2672
rect 294 2668 298 2672
rect 318 2668 322 2672
rect 342 2668 346 2672
rect 358 2668 362 2672
rect 374 2668 378 2672
rect 454 2668 458 2672
rect 558 2668 562 2672
rect 126 2658 130 2662
rect 198 2658 202 2662
rect 238 2658 242 2662
rect 246 2658 250 2662
rect 262 2658 266 2662
rect 302 2658 306 2662
rect 598 2668 602 2672
rect 710 2668 714 2672
rect 846 2668 850 2672
rect 854 2668 858 2672
rect 926 2668 930 2672
rect 942 2668 946 2672
rect 1054 2668 1058 2672
rect 1206 2668 1210 2672
rect 1238 2668 1242 2672
rect 1262 2668 1266 2672
rect 1334 2668 1338 2672
rect 1526 2668 1530 2672
rect 1646 2668 1650 2672
rect 1662 2668 1666 2672
rect 1734 2668 1738 2672
rect 1846 2668 1850 2672
rect 2062 2668 2066 2672
rect 2134 2668 2138 2672
rect 2230 2668 2234 2672
rect 2254 2668 2258 2672
rect 2270 2668 2274 2672
rect 2302 2668 2306 2672
rect 2318 2668 2322 2672
rect 2350 2668 2354 2672
rect 2366 2668 2370 2672
rect 2382 2668 2386 2672
rect 2406 2668 2410 2672
rect 2414 2668 2418 2672
rect 2462 2668 2466 2672
rect 2478 2668 2482 2672
rect 2598 2668 2602 2672
rect 2694 2668 2698 2672
rect 2726 2668 2730 2672
rect 2758 2668 2762 2672
rect 2766 2668 2770 2672
rect 2918 2668 2922 2672
rect 3006 2668 3010 2672
rect 3014 2668 3018 2672
rect 3022 2668 3026 2672
rect 3038 2668 3042 2672
rect 3070 2668 3074 2672
rect 3102 2668 3106 2672
rect 414 2658 418 2662
rect 462 2658 466 2662
rect 510 2658 514 2662
rect 550 2658 554 2662
rect 582 2658 586 2662
rect 590 2658 594 2662
rect 638 2658 642 2662
rect 766 2658 770 2662
rect 838 2658 842 2662
rect 862 2658 866 2662
rect 950 2658 954 2662
rect 998 2658 1002 2662
rect 1126 2658 1130 2662
rect 1150 2658 1154 2662
rect 1198 2658 1202 2662
rect 1286 2658 1290 2662
rect 1478 2658 1482 2662
rect 1582 2658 1586 2662
rect 1654 2658 1658 2662
rect 1694 2658 1698 2662
rect 1878 2658 1882 2662
rect 1910 2658 1914 2662
rect 2102 2658 2106 2662
rect 2142 2658 2146 2662
rect 2166 2658 2170 2662
rect 2174 2658 2178 2662
rect 2198 2658 2202 2662
rect 2206 2658 2210 2662
rect 2294 2658 2298 2662
rect 2310 2658 2314 2662
rect 2326 2658 2330 2662
rect 2342 2658 2346 2662
rect 2374 2658 2378 2662
rect 3134 2668 3138 2672
rect 3166 2668 3170 2672
rect 3182 2668 3186 2672
rect 3230 2668 3234 2672
rect 3246 2668 3250 2672
rect 3262 2668 3266 2672
rect 3286 2668 3290 2672
rect 3414 2668 3418 2672
rect 3534 2668 3538 2672
rect 3558 2668 3562 2672
rect 3574 2668 3578 2672
rect 3606 2668 3610 2672
rect 3678 2668 3682 2672
rect 3702 2668 3706 2672
rect 3710 2668 3714 2672
rect 3758 2668 3762 2672
rect 3782 2668 3786 2672
rect 3790 2668 3794 2672
rect 3814 2668 3818 2672
rect 3830 2668 3834 2672
rect 3862 2678 3866 2682
rect 3990 2678 3994 2682
rect 3998 2678 4002 2682
rect 4190 2678 4194 2682
rect 3886 2668 3890 2672
rect 3918 2668 3922 2672
rect 3934 2668 3938 2672
rect 4006 2668 4010 2672
rect 4038 2668 4042 2672
rect 4046 2668 4050 2672
rect 4094 2668 4098 2672
rect 4126 2668 4130 2672
rect 4182 2668 4186 2672
rect 4246 2668 4250 2672
rect 4254 2668 4258 2672
rect 2438 2658 2442 2662
rect 2470 2658 2474 2662
rect 2542 2658 2546 2662
rect 2670 2658 2674 2662
rect 2702 2658 2706 2662
rect 2718 2658 2722 2662
rect 2734 2658 2738 2662
rect 2750 2658 2754 2662
rect 2790 2658 2794 2662
rect 2950 2658 2954 2662
rect 3046 2658 3050 2662
rect 3062 2658 3066 2662
rect 3078 2658 3082 2662
rect 3094 2658 3098 2662
rect 3110 2658 3114 2662
rect 3126 2658 3130 2662
rect 3158 2658 3162 2662
rect 3174 2658 3178 2662
rect 3222 2658 3226 2662
rect 3238 2658 3242 2662
rect 3278 2658 3282 2662
rect 3310 2658 3314 2662
rect 3334 2658 3338 2662
rect 3342 2658 3346 2662
rect 3366 2658 3370 2662
rect 3518 2658 3522 2662
rect 3542 2658 3546 2662
rect 3566 2658 3570 2662
rect 3598 2658 3602 2662
rect 3614 2658 3618 2662
rect 3638 2658 3642 2662
rect 3662 2658 3666 2662
rect 3670 2658 3674 2662
rect 3710 2658 3714 2662
rect 3742 2658 3746 2662
rect 3750 2658 3754 2662
rect 3822 2658 3826 2662
rect 3894 2658 3898 2662
rect 4286 2668 4290 2672
rect 4334 2668 4338 2672
rect 4342 2668 4346 2672
rect 4390 2668 4394 2672
rect 3958 2658 3962 2662
rect 4014 2658 4018 2662
rect 4118 2658 4122 2662
rect 4142 2658 4146 2662
rect 4230 2658 4234 2662
rect 4262 2658 4266 2662
rect 4278 2658 4282 2662
rect 4302 2658 4306 2662
rect 38 2650 42 2654
rect 166 2648 170 2652
rect 246 2648 250 2652
rect 278 2648 282 2652
rect 526 2648 530 2652
rect 534 2648 538 2652
rect 566 2648 570 2652
rect 614 2648 618 2652
rect 678 2650 682 2654
rect 822 2648 826 2652
rect 878 2648 882 2652
rect 902 2648 906 2652
rect 1086 2650 1090 2654
rect 1182 2648 1186 2652
rect 1214 2648 1218 2652
rect 1246 2648 1250 2652
rect 1302 2650 1306 2654
rect 1494 2650 1498 2654
rect 1638 2648 1642 2652
rect 1702 2650 1706 2654
rect 1854 2648 1858 2652
rect 2094 2650 2098 2654
rect 2158 2648 2162 2652
rect 2214 2648 2218 2652
rect 2326 2648 2330 2652
rect 2358 2648 2362 2652
rect 2486 2648 2490 2652
rect 2630 2650 2634 2654
rect 2718 2648 2722 2652
rect 2806 2648 2810 2652
rect 2966 2648 2970 2652
rect 3062 2648 3066 2652
rect 3110 2648 3114 2652
rect 3142 2648 3146 2652
rect 3206 2648 3210 2652
rect 3294 2648 3298 2652
rect 3382 2650 3386 2654
rect 3582 2648 3586 2652
rect 3726 2648 3730 2652
rect 3766 2648 3770 2652
rect 3774 2648 3778 2652
rect 3806 2648 3810 2652
rect 3838 2648 3842 2652
rect 3910 2648 3914 2652
rect 3934 2648 3938 2652
rect 3966 2648 3970 2652
rect 4102 2648 4106 2652
rect 4134 2648 4138 2652
rect 4278 2648 4282 2652
rect 1838 2638 1842 2642
rect 1950 2638 1954 2642
rect 3518 2638 3522 2642
rect 3950 2638 3954 2642
rect 4150 2638 4154 2642
rect 4166 2638 4170 2642
rect 126 2627 130 2631
rect 766 2627 770 2631
rect 998 2627 1002 2631
rect 1302 2627 1306 2631
rect 1702 2627 1706 2631
rect 2278 2628 2282 2632
rect 2630 2627 2634 2631
rect 3958 2628 3962 2632
rect 510 2618 514 2622
rect 1430 2618 1434 2622
rect 1494 2618 1498 2622
rect 1894 2618 1898 2622
rect 2094 2618 2098 2622
rect 2238 2618 2242 2622
rect 2502 2618 2506 2622
rect 2822 2618 2826 2622
rect 2966 2618 2970 2622
rect 3326 2618 3330 2622
rect 3382 2618 3386 2622
rect 3694 2618 3698 2622
rect 3846 2618 3850 2622
rect 3894 2618 3898 2622
rect 4078 2618 4082 2622
rect 4142 2618 4146 2622
rect 4358 2618 4362 2622
rect 394 2603 398 2607
rect 401 2603 405 2607
rect 1418 2603 1422 2607
rect 1425 2603 1429 2607
rect 2442 2603 2446 2607
rect 2449 2603 2453 2607
rect 3474 2603 3478 2607
rect 3481 2603 3485 2607
rect 278 2588 282 2592
rect 486 2588 490 2592
rect 542 2588 546 2592
rect 566 2588 570 2592
rect 606 2588 610 2592
rect 646 2588 650 2592
rect 670 2588 674 2592
rect 822 2588 826 2592
rect 854 2588 858 2592
rect 1046 2588 1050 2592
rect 1542 2588 1546 2592
rect 1766 2588 1770 2592
rect 1846 2588 1850 2592
rect 2142 2588 2146 2592
rect 2270 2588 2274 2592
rect 2318 2588 2322 2592
rect 2430 2588 2434 2592
rect 2518 2588 2522 2592
rect 2638 2588 2642 2592
rect 2670 2588 2674 2592
rect 3014 2588 3018 2592
rect 3086 2588 3090 2592
rect 3110 2588 3114 2592
rect 3238 2588 3242 2592
rect 3510 2588 3514 2592
rect 3926 2588 3930 2592
rect 3950 2588 3954 2592
rect 374 2578 378 2582
rect 790 2578 794 2582
rect 918 2579 922 2583
rect 1270 2579 1274 2583
rect 1342 2579 1346 2583
rect 1622 2579 1626 2583
rect 2822 2579 2826 2583
rect 3886 2578 3890 2582
rect 518 2568 522 2572
rect 534 2568 538 2572
rect 1534 2568 1538 2572
rect 1806 2568 1810 2572
rect 1822 2568 1826 2572
rect 3142 2568 3146 2572
rect 4038 2568 4042 2572
rect 4054 2568 4058 2572
rect 110 2558 114 2562
rect 206 2558 210 2562
rect 238 2558 242 2562
rect 422 2558 426 2562
rect 550 2558 554 2562
rect 806 2558 810 2562
rect 838 2558 842 2562
rect 918 2556 922 2560
rect 1270 2556 1274 2560
rect 1342 2556 1346 2560
rect 1558 2558 1562 2562
rect 1622 2556 1626 2560
rect 2070 2558 2074 2562
rect 2086 2558 2090 2562
rect 2102 2558 2106 2562
rect 2158 2558 2162 2562
rect 2286 2558 2290 2562
rect 2334 2558 2338 2562
rect 2366 2558 2370 2562
rect 2414 2558 2418 2562
rect 2478 2558 2482 2562
rect 2502 2558 2506 2562
rect 2582 2558 2586 2562
rect 2654 2558 2658 2562
rect 2822 2556 2826 2560
rect 3014 2558 3018 2562
rect 3198 2558 3202 2562
rect 3254 2558 3258 2562
rect 3270 2558 3274 2562
rect 3310 2558 3314 2562
rect 3510 2558 3514 2562
rect 3686 2558 3690 2562
rect 3718 2558 3722 2562
rect 22 2548 26 2552
rect 94 2548 98 2552
rect 190 2548 194 2552
rect 198 2548 202 2552
rect 214 2548 218 2552
rect 254 2548 258 2552
rect 374 2548 378 2552
rect 518 2548 522 2552
rect 542 2548 546 2552
rect 590 2548 594 2552
rect 622 2548 626 2552
rect 822 2548 826 2552
rect 862 2548 866 2552
rect 1006 2548 1010 2552
rect 1102 2548 1106 2552
rect 1126 2548 1130 2552
rect 1286 2548 1290 2552
rect 1334 2548 1338 2552
rect 6 2538 10 2542
rect 30 2538 34 2542
rect 78 2538 82 2542
rect 1518 2548 1522 2552
rect 1542 2548 1546 2552
rect 1574 2548 1578 2552
rect 1606 2548 1610 2552
rect 1751 2548 1755 2552
rect 1830 2548 1834 2552
rect 1886 2548 1890 2552
rect 1894 2548 1898 2552
rect 1942 2548 1946 2552
rect 118 2538 122 2542
rect 126 2538 130 2542
rect 142 2538 146 2542
rect 158 2538 162 2542
rect 182 2538 186 2542
rect 262 2538 266 2542
rect 374 2538 378 2542
rect 494 2538 498 2542
rect 726 2538 730 2542
rect 830 2538 834 2542
rect 870 2538 874 2542
rect 950 2538 954 2542
rect 1078 2538 1082 2542
rect 1094 2538 1098 2542
rect 1110 2538 1114 2542
rect 1238 2538 1242 2542
rect 1374 2538 1378 2542
rect 1430 2538 1434 2542
rect 1502 2538 1506 2542
rect 1582 2538 1586 2542
rect 1654 2538 1658 2542
rect 1774 2538 1778 2542
rect 1782 2538 1786 2542
rect 1806 2538 1810 2542
rect 1918 2538 1922 2542
rect 2006 2548 2010 2552
rect 2030 2548 2034 2552
rect 2038 2548 2042 2552
rect 2054 2548 2058 2552
rect 2062 2548 2066 2552
rect 2086 2548 2090 2552
rect 2126 2548 2130 2552
rect 2142 2548 2146 2552
rect 2166 2548 2170 2552
rect 2198 2548 2202 2552
rect 2238 2548 2242 2552
rect 2278 2548 2282 2552
rect 2318 2548 2322 2552
rect 2350 2548 2354 2552
rect 2358 2548 2362 2552
rect 2438 2548 2442 2552
rect 2470 2548 2474 2552
rect 2510 2548 2514 2552
rect 2534 2548 2538 2552
rect 2550 2548 2554 2552
rect 2598 2548 2602 2552
rect 2606 2548 2610 2552
rect 2670 2548 2674 2552
rect 2838 2548 2842 2552
rect 2046 2538 2050 2542
rect 2078 2538 2082 2542
rect 2134 2538 2138 2542
rect 2174 2538 2178 2542
rect 2302 2538 2306 2542
rect 2310 2538 2314 2542
rect 2342 2538 2346 2542
rect 2398 2538 2402 2542
rect 2454 2538 2458 2542
rect 2486 2538 2490 2542
rect 2502 2538 2506 2542
rect 2510 2538 2514 2542
rect 2542 2538 2546 2542
rect 2558 2538 2562 2542
rect 3006 2548 3010 2552
rect 3070 2548 3074 2552
rect 3126 2548 3130 2552
rect 3142 2548 3146 2552
rect 3158 2548 3162 2552
rect 3190 2548 3194 2552
rect 3214 2548 3218 2552
rect 3230 2548 3234 2552
rect 3270 2548 3274 2552
rect 3278 2548 3282 2552
rect 3334 2548 3338 2552
rect 3342 2548 3346 2552
rect 3510 2548 3514 2552
rect 3582 2548 3586 2552
rect 3670 2548 3674 2552
rect 3710 2548 3714 2552
rect 3766 2548 3770 2552
rect 3790 2558 3794 2562
rect 3894 2558 3898 2562
rect 3966 2558 3970 2562
rect 4022 2558 4026 2562
rect 4070 2558 4074 2562
rect 4158 2558 4162 2562
rect 3814 2548 3818 2552
rect 2686 2538 2690 2542
rect 2790 2538 2794 2542
rect 2910 2538 2914 2542
rect 2966 2538 2970 2542
rect 3054 2538 3058 2542
rect 3102 2538 3106 2542
rect 3134 2538 3138 2542
rect 3182 2538 3186 2542
rect 3206 2538 3210 2542
rect 3230 2538 3234 2542
rect 3278 2538 3282 2542
rect 3286 2538 3290 2542
rect 3310 2538 3314 2542
rect 3318 2538 3322 2542
rect 3350 2538 3354 2542
rect 3462 2538 3466 2542
rect 3614 2538 3618 2542
rect 3630 2538 3634 2542
rect 3638 2538 3642 2542
rect 3662 2538 3666 2542
rect 3678 2538 3682 2542
rect 3718 2538 3722 2542
rect 3742 2538 3746 2542
rect 3758 2538 3762 2542
rect 3774 2538 3778 2542
rect 3806 2538 3810 2542
rect 3838 2538 3842 2542
rect 3910 2548 3914 2552
rect 3950 2548 3954 2552
rect 3966 2548 3970 2552
rect 4014 2548 4018 2552
rect 4030 2548 4034 2552
rect 4126 2548 4130 2552
rect 4198 2558 4202 2562
rect 4350 2558 4354 2562
rect 4374 2558 4378 2562
rect 4174 2548 4178 2552
rect 4238 2548 4242 2552
rect 4246 2548 4250 2552
rect 4342 2548 4346 2552
rect 3870 2538 3874 2542
rect 3942 2538 3946 2542
rect 4006 2538 4010 2542
rect 4054 2538 4058 2542
rect 4062 2538 4066 2542
rect 4078 2538 4082 2542
rect 4126 2538 4130 2542
rect 4134 2538 4138 2542
rect 4190 2538 4194 2542
rect 4214 2538 4218 2542
rect 4270 2538 4274 2542
rect 4318 2538 4322 2542
rect 4374 2538 4378 2542
rect 4390 2538 4394 2542
rect 174 2528 178 2532
rect 214 2528 218 2532
rect 230 2528 234 2532
rect 358 2528 362 2532
rect 502 2528 506 2532
rect 558 2528 562 2532
rect 574 2528 578 2532
rect 638 2528 642 2532
rect 654 2528 658 2532
rect 966 2528 970 2532
rect 1222 2528 1226 2532
rect 1390 2528 1394 2532
rect 1486 2528 1490 2532
rect 1670 2528 1674 2532
rect 1870 2528 1874 2532
rect 1974 2528 1978 2532
rect 1990 2528 1994 2532
rect 2022 2528 2026 2532
rect 2110 2528 2114 2532
rect 2214 2528 2218 2532
rect 2254 2528 2258 2532
rect 2262 2528 2266 2532
rect 2390 2528 2394 2532
rect 2422 2528 2426 2532
rect 2614 2528 2618 2532
rect 2646 2528 2650 2532
rect 2774 2528 2778 2532
rect 2862 2528 2866 2532
rect 2950 2528 2954 2532
rect 3158 2528 3162 2532
rect 3166 2528 3170 2532
rect 3246 2528 3250 2532
rect 3446 2528 3450 2532
rect 3598 2528 3602 2532
rect 3614 2528 3618 2532
rect 3654 2528 3658 2532
rect 3750 2528 3754 2532
rect 3830 2528 3834 2532
rect 3838 2528 3842 2532
rect 3862 2528 3866 2532
rect 3934 2528 3938 2532
rect 3990 2528 3994 2532
rect 4222 2528 4226 2532
rect 110 2518 114 2522
rect 238 2518 242 2522
rect 486 2518 490 2522
rect 670 2518 674 2522
rect 790 2518 794 2522
rect 1142 2518 1146 2522
rect 1518 2518 1522 2522
rect 1790 2518 1794 2522
rect 1814 2518 1818 2522
rect 1958 2518 1962 2522
rect 2118 2518 2122 2522
rect 2246 2518 2250 2522
rect 2294 2518 2298 2522
rect 2382 2518 2386 2522
rect 2414 2518 2418 2522
rect 2566 2518 2570 2522
rect 2694 2518 2698 2522
rect 3062 2518 3066 2522
rect 3366 2518 3370 2522
rect 3574 2518 3578 2522
rect 3622 2518 3626 2522
rect 3694 2518 3698 2522
rect 3822 2518 3826 2522
rect 3894 2518 3898 2522
rect 4102 2518 4106 2522
rect 4206 2518 4210 2522
rect 4230 2518 4234 2522
rect 4302 2518 4306 2522
rect 4358 2518 4362 2522
rect 4374 2518 4378 2522
rect 898 2503 902 2507
rect 905 2503 909 2507
rect 1930 2503 1934 2507
rect 1937 2503 1941 2507
rect 2954 2503 2958 2507
rect 2961 2503 2965 2507
rect 3978 2503 3982 2507
rect 3985 2503 3989 2507
rect 166 2488 170 2492
rect 190 2488 194 2492
rect 214 2488 218 2492
rect 390 2488 394 2492
rect 486 2488 490 2492
rect 566 2488 570 2492
rect 590 2488 594 2492
rect 606 2488 610 2492
rect 646 2488 650 2492
rect 1294 2488 1298 2492
rect 1382 2488 1386 2492
rect 1454 2488 1458 2492
rect 1534 2488 1538 2492
rect 1630 2488 1634 2492
rect 1662 2488 1666 2492
rect 1870 2488 1874 2492
rect 2174 2488 2178 2492
rect 2190 2488 2194 2492
rect 2230 2488 2234 2492
rect 2350 2488 2354 2492
rect 2366 2488 2370 2492
rect 2622 2488 2626 2492
rect 2694 2488 2698 2492
rect 2710 2488 2714 2492
rect 2830 2488 2834 2492
rect 3246 2488 3250 2492
rect 3286 2488 3290 2492
rect 3310 2488 3314 2492
rect 3358 2488 3362 2492
rect 3550 2488 3554 2492
rect 3718 2488 3722 2492
rect 3854 2488 3858 2492
rect 3886 2488 3890 2492
rect 4014 2488 4018 2492
rect 4190 2488 4194 2492
rect 4318 2488 4322 2492
rect 86 2478 90 2482
rect 294 2478 298 2482
rect 382 2478 386 2482
rect 494 2478 498 2482
rect 558 2478 562 2482
rect 582 2478 586 2482
rect 726 2478 730 2482
rect 926 2478 930 2482
rect 1046 2478 1050 2482
rect 1150 2478 1154 2482
rect 1334 2478 1338 2482
rect 1462 2478 1466 2482
rect 1726 2478 1730 2482
rect 1734 2478 1738 2482
rect 1766 2478 1770 2482
rect 2030 2478 2034 2482
rect 2038 2478 2042 2482
rect 2158 2478 2162 2482
rect 2166 2478 2170 2482
rect 2262 2478 2266 2482
rect 2406 2478 2410 2482
rect 2486 2478 2490 2482
rect 2582 2478 2586 2482
rect 3078 2478 3082 2482
rect 3086 2478 3090 2482
rect 3158 2478 3162 2482
rect 3182 2478 3186 2482
rect 3270 2478 3274 2482
rect 3278 2478 3282 2482
rect 3302 2478 3306 2482
rect 3422 2478 3426 2482
rect 3454 2478 3458 2482
rect 3502 2478 3506 2482
rect 3606 2478 3610 2482
rect 3662 2478 3666 2482
rect 3702 2478 3706 2482
rect 3782 2478 3786 2482
rect 3838 2478 3842 2482
rect 3966 2478 3970 2482
rect 4358 2478 4362 2482
rect 70 2468 74 2472
rect 310 2468 314 2472
rect 478 2468 482 2472
rect 502 2468 506 2472
rect 550 2468 554 2472
rect 630 2468 634 2472
rect 742 2468 746 2472
rect 814 2468 818 2472
rect 910 2468 914 2472
rect 1007 2468 1011 2472
rect 1134 2468 1138 2472
rect 1270 2468 1274 2472
rect 1374 2468 1378 2472
rect 1406 2468 1410 2472
rect 1470 2468 1474 2472
rect 1486 2468 1490 2472
rect 1526 2468 1530 2472
rect 1622 2468 1626 2472
rect 1654 2468 1658 2472
rect 1678 2468 1682 2472
rect 1686 2468 1690 2472
rect 1702 2468 1706 2472
rect 1718 2468 1722 2472
rect 1742 2468 1746 2472
rect 1798 2468 1802 2472
rect 1830 2468 1834 2472
rect 1942 2468 1946 2472
rect 1974 2468 1978 2472
rect 2006 2468 2010 2472
rect 2062 2468 2066 2472
rect 2078 2468 2082 2472
rect 2094 2468 2098 2472
rect 2102 2468 2106 2472
rect 2326 2468 2330 2472
rect 2374 2468 2378 2472
rect 2502 2468 2506 2472
rect 2598 2468 2602 2472
rect 2614 2468 2618 2472
rect 2646 2468 2650 2472
rect 2654 2468 2658 2472
rect 2686 2468 2690 2472
rect 2702 2468 2706 2472
rect 2718 2468 2722 2472
rect 2734 2468 2738 2472
rect 2750 2468 2754 2472
rect 2774 2468 2778 2472
rect 2806 2468 2810 2472
rect 2894 2468 2898 2472
rect 2910 2468 2914 2472
rect 2926 2468 2930 2472
rect 3038 2468 3042 2472
rect 3094 2468 3098 2472
rect 3110 2468 3114 2472
rect 3126 2468 3130 2472
rect 3166 2468 3170 2472
rect 3214 2468 3218 2472
rect 3222 2468 3226 2472
rect 126 2458 130 2462
rect 254 2458 258 2462
rect 406 2458 410 2462
rect 542 2458 546 2462
rect 574 2458 578 2462
rect 622 2458 626 2462
rect 782 2458 786 2462
rect 966 2458 970 2462
rect 1062 2458 1066 2462
rect 1086 2458 1090 2462
rect 1238 2458 1242 2462
rect 1278 2458 1282 2462
rect 1318 2458 1322 2462
rect 1350 2458 1354 2462
rect 1366 2458 1370 2462
rect 1398 2458 1402 2462
rect 1430 2458 1434 2462
rect 1438 2458 1442 2462
rect 1502 2458 1506 2462
rect 1582 2458 1586 2462
rect 1614 2458 1618 2462
rect 1646 2458 1650 2462
rect 1694 2458 1698 2462
rect 1710 2458 1714 2462
rect 1750 2458 1754 2462
rect 1822 2458 1826 2462
rect 1854 2458 1858 2462
rect 1894 2458 1898 2462
rect 1918 2458 1922 2462
rect 1950 2458 1954 2462
rect 1966 2458 1970 2462
rect 1982 2458 1986 2462
rect 1998 2458 2002 2462
rect 2014 2458 2018 2462
rect 2022 2458 2026 2462
rect 2054 2458 2058 2462
rect 2086 2458 2090 2462
rect 2110 2458 2114 2462
rect 2126 2458 2130 2462
rect 2142 2458 2146 2462
rect 2214 2458 2218 2462
rect 2222 2458 2226 2462
rect 2246 2458 2250 2462
rect 2254 2458 2258 2462
rect 2262 2458 2266 2462
rect 2310 2458 2314 2462
rect 2318 2458 2322 2462
rect 2334 2458 2338 2462
rect 2446 2458 2450 2462
rect 2534 2458 2538 2462
rect 2606 2458 2610 2462
rect 2638 2458 2642 2462
rect 2662 2458 2666 2462
rect 2678 2458 2682 2462
rect 2726 2458 2730 2462
rect 2774 2458 2778 2462
rect 2782 2458 2786 2462
rect 2814 2458 2818 2462
rect 2846 2458 2850 2462
rect 2854 2458 2858 2462
rect 2878 2458 2882 2462
rect 2902 2458 2906 2462
rect 2918 2458 2922 2462
rect 2950 2458 2954 2462
rect 2958 2458 2962 2462
rect 2982 2458 2986 2462
rect 2998 2458 3002 2462
rect 3006 2458 3010 2462
rect 3030 2458 3034 2462
rect 3070 2458 3074 2462
rect 3374 2468 3378 2472
rect 3414 2468 3418 2472
rect 3438 2468 3442 2472
rect 3526 2468 3530 2472
rect 3630 2468 3634 2472
rect 3646 2468 3650 2472
rect 3694 2468 3698 2472
rect 3710 2468 3714 2472
rect 3774 2468 3778 2472
rect 3846 2468 3850 2472
rect 3870 2468 3874 2472
rect 3918 2468 3922 2472
rect 3982 2468 3986 2472
rect 4022 2468 4026 2472
rect 4078 2468 4082 2472
rect 4134 2468 4138 2472
rect 4150 2468 4154 2472
rect 4198 2468 4202 2472
rect 4230 2468 4234 2472
rect 4238 2468 4242 2472
rect 4334 2468 4338 2472
rect 4390 2468 4394 2472
rect 3118 2458 3122 2462
rect 3142 2458 3146 2462
rect 3166 2458 3170 2462
rect 3206 2458 3210 2462
rect 3214 2458 3218 2462
rect 3254 2458 3258 2462
rect 3294 2458 3298 2462
rect 3318 2458 3322 2462
rect 3350 2458 3354 2462
rect 3366 2458 3370 2462
rect 3398 2458 3402 2462
rect 3414 2458 3418 2462
rect 3446 2458 3450 2462
rect 3486 2458 3490 2462
rect 3494 2458 3498 2462
rect 3518 2458 3522 2462
rect 3534 2458 3538 2462
rect 3558 2458 3562 2462
rect 3566 2458 3570 2462
rect 3590 2458 3594 2462
rect 3622 2458 3626 2462
rect 3638 2458 3642 2462
rect 3670 2458 3674 2462
rect 3726 2458 3730 2462
rect 3766 2458 3770 2462
rect 3814 2458 3818 2462
rect 3926 2458 3930 2462
rect 3950 2458 3954 2462
rect 4078 2458 4082 2462
rect 4118 2458 4122 2462
rect 4158 2458 4162 2462
rect 4222 2458 4226 2462
rect 4286 2458 4290 2462
rect 4342 2458 4346 2462
rect 4358 2458 4362 2462
rect 4374 2458 4378 2462
rect 4382 2458 4386 2462
rect 38 2450 42 2454
rect 358 2448 362 2452
rect 502 2448 506 2452
rect 526 2448 530 2452
rect 606 2448 610 2452
rect 774 2450 778 2454
rect 878 2450 882 2454
rect 1102 2450 1106 2454
rect 1326 2448 1330 2452
rect 1350 2448 1354 2452
rect 1382 2448 1386 2452
rect 1454 2448 1458 2452
rect 1494 2448 1498 2452
rect 1598 2448 1602 2452
rect 1630 2448 1634 2452
rect 1662 2448 1666 2452
rect 1774 2448 1778 2452
rect 1966 2448 1970 2452
rect 2038 2448 2042 2452
rect 2070 2448 2074 2452
rect 2350 2448 2354 2452
rect 2358 2448 2362 2452
rect 2550 2448 2554 2452
rect 2590 2448 2594 2452
rect 2622 2448 2626 2452
rect 2742 2448 2746 2452
rect 2750 2448 2754 2452
rect 3134 2448 3138 2452
rect 3190 2448 3194 2452
rect 3206 2448 3210 2452
rect 3246 2448 3250 2452
rect 3334 2448 3338 2452
rect 3470 2448 3474 2452
rect 3550 2448 3554 2452
rect 3606 2448 3610 2452
rect 3798 2448 3802 2452
rect 4014 2448 4018 2452
rect 4070 2448 4074 2452
rect 4174 2448 4178 2452
rect 4182 2448 4186 2452
rect 4206 2448 4210 2452
rect 4270 2448 4274 2452
rect 4318 2448 4322 2452
rect 4366 2448 4370 2452
rect 1310 2438 1314 2442
rect 1510 2438 1514 2442
rect 1550 2438 1554 2442
rect 1574 2438 1578 2442
rect 3254 2438 3258 2442
rect 4158 2438 4162 2442
rect 126 2427 130 2431
rect 254 2427 258 2431
rect 774 2427 778 2431
rect 878 2427 882 2431
rect 1102 2427 1106 2431
rect 1582 2428 1586 2432
rect 3142 2428 3146 2432
rect 3662 2428 3666 2432
rect 822 2418 826 2422
rect 1030 2418 1034 2422
rect 1230 2418 1234 2422
rect 1342 2418 1346 2422
rect 1478 2418 1482 2422
rect 1502 2418 1506 2422
rect 1758 2418 1762 2422
rect 1782 2418 1786 2422
rect 1806 2418 1810 2422
rect 1910 2418 1914 2422
rect 1990 2418 1994 2422
rect 2118 2418 2122 2422
rect 2302 2418 2306 2422
rect 2550 2418 2554 2422
rect 2574 2418 2578 2422
rect 2870 2418 2874 2422
rect 2974 2418 2978 2422
rect 3022 2418 3026 2422
rect 3406 2418 3410 2422
rect 3582 2418 3586 2422
rect 3830 2418 3834 2422
rect 3902 2418 3906 2422
rect 4046 2418 4050 2422
rect 4102 2418 4106 2422
rect 4222 2418 4226 2422
rect 4246 2418 4250 2422
rect 394 2403 398 2407
rect 401 2403 405 2407
rect 1418 2403 1422 2407
rect 1425 2403 1429 2407
rect 2442 2403 2446 2407
rect 2449 2403 2453 2407
rect 3474 2403 3478 2407
rect 3481 2403 3485 2407
rect 182 2388 186 2392
rect 438 2388 442 2392
rect 478 2388 482 2392
rect 646 2388 650 2392
rect 1054 2388 1058 2392
rect 1182 2388 1186 2392
rect 1350 2388 1354 2392
rect 1638 2388 1642 2392
rect 1742 2388 1746 2392
rect 1798 2388 1802 2392
rect 1830 2388 1834 2392
rect 1982 2388 1986 2392
rect 2014 2388 2018 2392
rect 2486 2388 2490 2392
rect 2718 2388 2722 2392
rect 2750 2388 2754 2392
rect 2854 2388 2858 2392
rect 2934 2388 2938 2392
rect 3142 2388 3146 2392
rect 3638 2388 3642 2392
rect 4294 2388 4298 2392
rect 310 2379 314 2383
rect 518 2379 522 2383
rect 814 2379 818 2383
rect 902 2379 906 2383
rect 1222 2379 1226 2383
rect 2390 2379 2394 2383
rect 3502 2379 3506 2383
rect 1086 2368 1090 2372
rect 1126 2368 1130 2372
rect 1174 2368 1178 2372
rect 1438 2368 1442 2372
rect 1454 2368 1458 2372
rect 1654 2368 1658 2372
rect 1790 2368 1794 2372
rect 2590 2368 2594 2372
rect 2638 2368 2642 2372
rect 2806 2368 2810 2372
rect 3182 2368 3186 2372
rect 182 2358 186 2362
rect 310 2356 314 2360
rect 518 2356 522 2360
rect 814 2356 818 2360
rect 878 2358 882 2362
rect 6 2348 10 2352
rect 22 2348 26 2352
rect 182 2348 186 2352
rect 294 2348 298 2352
rect 606 2348 610 2352
rect 782 2348 786 2352
rect 830 2348 834 2352
rect 902 2356 906 2360
rect 1102 2358 1106 2362
rect 1110 2358 1114 2362
rect 1158 2358 1162 2362
rect 1222 2356 1226 2360
rect 1358 2358 1362 2362
rect 1694 2358 1698 2362
rect 1782 2358 1786 2362
rect 1806 2358 1810 2362
rect 2006 2358 2010 2362
rect 2070 2358 2074 2362
rect 2126 2358 2130 2362
rect 2158 2358 2162 2362
rect 2238 2358 2242 2362
rect 2390 2356 2394 2360
rect 2470 2358 2474 2362
rect 990 2348 994 2352
rect 1054 2348 1058 2352
rect 1094 2348 1098 2352
rect 1126 2348 1130 2352
rect 1166 2348 1170 2352
rect 1214 2348 1218 2352
rect 1374 2348 1378 2352
rect 1382 2348 1386 2352
rect 1470 2348 1474 2352
rect 1486 2348 1490 2352
rect 1526 2348 1530 2352
rect 1542 2348 1546 2352
rect 1646 2348 1650 2352
rect 1654 2348 1658 2352
rect 1670 2348 1674 2352
rect 1710 2348 1714 2352
rect 1726 2348 1730 2352
rect 1750 2348 1754 2352
rect 1782 2348 1786 2352
rect 1814 2348 1818 2352
rect 1846 2348 1850 2352
rect 1878 2348 1882 2352
rect 1886 2348 1890 2352
rect 1934 2348 1938 2352
rect 1950 2348 1954 2352
rect 1974 2348 1978 2352
rect 1998 2348 2002 2352
rect 2030 2348 2034 2352
rect 2070 2348 2074 2352
rect 2086 2348 2090 2352
rect 2110 2348 2114 2352
rect 2134 2348 2138 2352
rect 2142 2348 2146 2352
rect 2174 2348 2178 2352
rect 2190 2348 2194 2352
rect 2206 2348 2210 2352
rect 2230 2348 2234 2352
rect 2406 2348 2410 2352
rect 2454 2348 2458 2352
rect 2470 2348 2474 2352
rect 2502 2358 2506 2362
rect 2518 2348 2522 2352
rect 2526 2348 2530 2352
rect 2542 2348 2546 2352
rect 2566 2358 2570 2362
rect 2606 2358 2610 2362
rect 2654 2358 2658 2362
rect 2662 2358 2666 2362
rect 2790 2358 2794 2362
rect 2838 2358 2842 2362
rect 2870 2358 2874 2362
rect 2902 2358 2906 2362
rect 2998 2358 3002 2362
rect 3054 2358 3058 2362
rect 3166 2358 3170 2362
rect 2638 2348 2642 2352
rect 2678 2348 2682 2352
rect 2734 2348 2738 2352
rect 2774 2348 2778 2352
rect 2790 2348 2794 2352
rect 2822 2348 2826 2352
rect 2838 2348 2842 2352
rect 2854 2348 2858 2352
rect 2886 2348 2890 2352
rect 3502 2356 3506 2360
rect 3550 2358 3554 2362
rect 3574 2358 3578 2362
rect 3638 2358 3642 2362
rect 3814 2358 3818 2362
rect 3838 2358 3842 2362
rect 3894 2358 3898 2362
rect 4054 2358 4058 2362
rect 2934 2348 2938 2352
rect 2990 2348 2994 2352
rect 3014 2348 3018 2352
rect 3022 2348 3026 2352
rect 3046 2348 3050 2352
rect 3054 2348 3058 2352
rect 3070 2348 3074 2352
rect 3086 2348 3090 2352
rect 3094 2348 3098 2352
rect 3118 2348 3122 2352
rect 3158 2348 3162 2352
rect 3182 2348 3186 2352
rect 3198 2348 3202 2352
rect 3230 2348 3234 2352
rect 3254 2348 3258 2352
rect 3262 2348 3266 2352
rect 3294 2348 3298 2352
rect 3302 2348 3306 2352
rect 3350 2348 3354 2352
rect 3414 2348 3418 2352
rect 3510 2348 3514 2352
rect 3518 2348 3522 2352
rect 3574 2348 3578 2352
rect 3590 2348 3594 2352
rect 3638 2348 3642 2352
rect 3838 2348 3842 2352
rect 3902 2348 3906 2352
rect 3998 2348 4002 2352
rect 4046 2348 4050 2352
rect 4102 2358 4106 2362
rect 4150 2358 4154 2362
rect 4182 2358 4186 2362
rect 4198 2358 4202 2362
rect 4134 2348 4138 2352
rect 4182 2348 4186 2352
rect 4214 2348 4218 2352
rect 4238 2358 4242 2362
rect 4286 2358 4290 2362
rect 4390 2358 4394 2362
rect 4262 2348 4266 2352
rect 4310 2348 4314 2352
rect 4342 2348 4346 2352
rect 4374 2348 4378 2352
rect 22 2338 26 2342
rect 134 2338 138 2342
rect 206 2338 210 2342
rect 342 2338 346 2342
rect 550 2338 554 2342
rect 726 2338 730 2342
rect 782 2338 786 2342
rect 934 2338 938 2342
rect 1046 2338 1050 2342
rect 1134 2338 1138 2342
rect 1150 2338 1154 2342
rect 1254 2338 1258 2342
rect 1390 2338 1394 2342
rect 1398 2338 1402 2342
rect 1438 2338 1442 2342
rect 1462 2338 1466 2342
rect 1478 2338 1482 2342
rect 1494 2338 1498 2342
rect 1518 2338 1522 2342
rect 1550 2338 1554 2342
rect 1646 2338 1650 2342
rect 1678 2338 1682 2342
rect 1702 2338 1706 2342
rect 1734 2338 1738 2342
rect 1766 2338 1770 2342
rect 1822 2338 1826 2342
rect 1854 2338 1858 2342
rect 1870 2338 1874 2342
rect 1910 2338 1914 2342
rect 1966 2338 1970 2342
rect 2022 2338 2026 2342
rect 2030 2338 2034 2342
rect 2062 2338 2066 2342
rect 2078 2338 2082 2342
rect 2102 2338 2106 2342
rect 2134 2338 2138 2342
rect 2182 2338 2186 2342
rect 2358 2338 2362 2342
rect 2446 2338 2450 2342
rect 2478 2338 2482 2342
rect 2534 2338 2538 2342
rect 2582 2338 2586 2342
rect 2590 2338 2594 2342
rect 2630 2338 2634 2342
rect 2686 2338 2690 2342
rect 2694 2338 2698 2342
rect 2758 2338 2762 2342
rect 2766 2338 2770 2342
rect 2798 2338 2802 2342
rect 2846 2338 2850 2342
rect 2878 2338 2882 2342
rect 2902 2338 2906 2342
rect 2910 2338 2914 2342
rect 2982 2338 2986 2342
rect 3078 2338 3082 2342
rect 3126 2338 3130 2342
rect 3190 2338 3194 2342
rect 3206 2338 3210 2342
rect 3238 2338 3242 2342
rect 3270 2338 3274 2342
rect 3286 2338 3290 2342
rect 3310 2338 3314 2342
rect 3326 2338 3330 2342
rect 3358 2338 3362 2342
rect 3470 2338 3474 2342
rect 3582 2338 3586 2342
rect 3598 2338 3602 2342
rect 3686 2338 3690 2342
rect 3798 2338 3802 2342
rect 3822 2338 3826 2342
rect 3870 2338 3874 2342
rect 3894 2338 3898 2342
rect 3926 2338 3930 2342
rect 4014 2338 4018 2342
rect 4070 2338 4074 2342
rect 4118 2338 4122 2342
rect 4206 2338 4210 2342
rect 4222 2338 4226 2342
rect 4254 2338 4258 2342
rect 4302 2338 4306 2342
rect 4334 2338 4338 2342
rect 4358 2338 4362 2342
rect 4382 2338 4386 2342
rect 118 2328 122 2332
rect 358 2328 362 2332
rect 470 2328 474 2332
rect 566 2328 570 2332
rect 766 2328 770 2332
rect 950 2328 954 2332
rect 1270 2328 1274 2332
rect 1502 2328 1506 2332
rect 1542 2328 1546 2332
rect 1622 2328 1626 2332
rect 1694 2328 1698 2332
rect 1750 2328 1754 2332
rect 1838 2328 1842 2332
rect 2222 2328 2226 2332
rect 2246 2328 2250 2332
rect 2342 2328 2346 2332
rect 2558 2328 2562 2332
rect 2614 2328 2618 2332
rect 2702 2328 2706 2332
rect 2966 2328 2970 2332
rect 2998 2328 3002 2332
rect 3030 2328 3034 2332
rect 3222 2328 3226 2332
rect 3286 2328 3290 2332
rect 3326 2328 3330 2332
rect 3454 2328 3458 2332
rect 3614 2328 3618 2332
rect 3702 2328 3706 2332
rect 3862 2328 3866 2332
rect 4014 2328 4018 2332
rect 4158 2328 4162 2332
rect 262 2318 266 2322
rect 670 2318 674 2322
rect 686 2318 690 2322
rect 1030 2318 1034 2322
rect 1406 2318 1410 2322
rect 1446 2318 1450 2322
rect 1510 2318 1514 2322
rect 1606 2318 1610 2322
rect 1726 2318 1730 2322
rect 1862 2318 1866 2322
rect 1902 2318 1906 2322
rect 2046 2318 2050 2322
rect 2262 2318 2266 2322
rect 2662 2318 2666 2322
rect 2750 2318 2754 2322
rect 3214 2318 3218 2322
rect 3374 2318 3378 2322
rect 3606 2318 3610 2322
rect 3782 2318 3786 2322
rect 3814 2318 3818 2322
rect 3830 2318 3834 2322
rect 3854 2318 3858 2322
rect 3886 2318 3890 2322
rect 3918 2318 3922 2322
rect 3958 2318 3962 2322
rect 4086 2318 4090 2322
rect 4150 2318 4154 2322
rect 4350 2318 4354 2322
rect 898 2303 902 2307
rect 905 2303 909 2307
rect 1930 2303 1934 2307
rect 1937 2303 1941 2307
rect 2954 2303 2958 2307
rect 2961 2303 2965 2307
rect 3978 2303 3982 2307
rect 3985 2303 3989 2307
rect 6 2288 10 2292
rect 62 2288 66 2292
rect 750 2288 754 2292
rect 782 2288 786 2292
rect 886 2288 890 2292
rect 1006 2288 1010 2292
rect 1038 2288 1042 2292
rect 1062 2288 1066 2292
rect 1094 2288 1098 2292
rect 1318 2288 1322 2292
rect 1334 2288 1338 2292
rect 1582 2288 1586 2292
rect 1638 2288 1642 2292
rect 1710 2288 1714 2292
rect 2022 2288 2026 2292
rect 2326 2288 2330 2292
rect 2454 2288 2458 2292
rect 2830 2288 2834 2292
rect 3342 2288 3346 2292
rect 3590 2288 3594 2292
rect 3686 2288 3690 2292
rect 4190 2288 4194 2292
rect 174 2278 178 2282
rect 350 2278 354 2282
rect 534 2278 538 2282
rect 1014 2278 1018 2282
rect 1206 2278 1210 2282
rect 1454 2278 1458 2282
rect 1550 2278 1554 2282
rect 1614 2278 1618 2282
rect 1622 2278 1626 2282
rect 1718 2278 1722 2282
rect 1814 2278 1818 2282
rect 1854 2278 1858 2282
rect 1878 2278 1882 2282
rect 1990 2278 1994 2282
rect 2038 2278 2042 2282
rect 2094 2278 2098 2282
rect 2118 2278 2122 2282
rect 2214 2278 2218 2282
rect 2334 2278 2338 2282
rect 2390 2278 2394 2282
rect 2406 2278 2410 2282
rect 2550 2278 2554 2282
rect 2734 2278 2738 2282
rect 2926 2278 2930 2282
rect 3118 2278 3122 2282
rect 3422 2278 3426 2282
rect 3502 2278 3506 2282
rect 3614 2278 3618 2282
rect 3918 2278 3922 2282
rect 3990 2278 3994 2282
rect 4006 2278 4010 2282
rect 4182 2278 4186 2282
rect 4198 2278 4202 2282
rect 4254 2278 4258 2282
rect 4294 2278 4298 2282
rect 4310 2278 4314 2282
rect 4350 2278 4354 2282
rect 22 2268 26 2272
rect 190 2268 194 2272
rect 366 2268 370 2272
rect 518 2268 522 2272
rect 622 2268 626 2272
rect 646 2268 650 2272
rect 662 2268 666 2272
rect 678 2268 682 2272
rect 694 2268 698 2272
rect 710 2268 714 2272
rect 726 2268 730 2272
rect 758 2268 762 2272
rect 822 2268 826 2272
rect 910 2268 914 2272
rect 926 2268 930 2272
rect 958 2268 962 2272
rect 974 2268 978 2272
rect 982 2268 986 2272
rect 1054 2268 1058 2272
rect 1086 2268 1090 2272
rect 1118 2268 1122 2272
rect 1190 2268 1194 2272
rect 1302 2268 1306 2272
rect 1438 2268 1442 2272
rect 1590 2268 1594 2272
rect 1606 2268 1610 2272
rect 1630 2268 1634 2272
rect 1662 2268 1666 2272
rect 1670 2268 1674 2272
rect 1702 2268 1706 2272
rect 1726 2268 1730 2272
rect 1774 2268 1778 2272
rect 1814 2268 1818 2272
rect 1886 2268 1890 2272
rect 1918 2268 1922 2272
rect 1966 2268 1970 2272
rect 1990 2268 1994 2272
rect 2038 2268 2042 2272
rect 2230 2268 2234 2272
rect 2302 2268 2306 2272
rect 2414 2268 2418 2272
rect 2454 2268 2458 2272
rect 2494 2268 2498 2272
rect 2526 2268 2530 2272
rect 2550 2268 2554 2272
rect 2590 2268 2594 2272
rect 2750 2268 2754 2272
rect 2822 2268 2826 2272
rect 2886 2268 2890 2272
rect 2942 2268 2946 2272
rect 3078 2268 3082 2272
rect 3134 2268 3138 2272
rect 3214 2268 3218 2272
rect 3230 2268 3234 2272
rect 3246 2268 3250 2272
rect 3302 2268 3306 2272
rect 3318 2268 3322 2272
rect 3334 2268 3338 2272
rect 3390 2268 3394 2272
rect 3406 2268 3410 2272
rect 3454 2268 3458 2272
rect 3486 2268 3490 2272
rect 3534 2268 3538 2272
rect 3566 2268 3570 2272
rect 3582 2268 3586 2272
rect 3606 2268 3610 2272
rect 3630 2268 3634 2272
rect 3670 2268 3674 2272
rect 3678 2268 3682 2272
rect 3702 2268 3706 2272
rect 3718 2268 3722 2272
rect 3742 2268 3746 2272
rect 3822 2268 3826 2272
rect 3862 2268 3866 2272
rect 3942 2268 3946 2272
rect 4014 2268 4018 2272
rect 4030 2268 4034 2272
rect 4094 2268 4098 2272
rect 4142 2268 4146 2272
rect 4158 2268 4162 2272
rect 4174 2268 4178 2272
rect 4214 2268 4218 2272
rect 4222 2268 4226 2272
rect 4286 2268 4290 2272
rect 4342 2268 4346 2272
rect 4366 2268 4370 2272
rect 38 2258 42 2262
rect 222 2258 226 2262
rect 414 2258 418 2262
rect 6 2248 10 2252
rect 22 2248 26 2252
rect 238 2248 242 2252
rect 398 2250 402 2254
rect 574 2258 578 2262
rect 670 2258 674 2262
rect 726 2258 730 2262
rect 734 2258 738 2262
rect 766 2258 770 2262
rect 806 2258 810 2262
rect 830 2258 834 2262
rect 846 2258 850 2262
rect 870 2258 874 2262
rect 902 2258 906 2262
rect 950 2258 954 2262
rect 1030 2258 1034 2262
rect 1078 2258 1082 2262
rect 1110 2258 1114 2262
rect 1246 2258 1250 2262
rect 1342 2258 1346 2262
rect 1390 2258 1394 2262
rect 1494 2258 1498 2262
rect 1566 2258 1570 2262
rect 1598 2258 1602 2262
rect 1638 2258 1642 2262
rect 1662 2258 1666 2262
rect 1678 2258 1682 2262
rect 1694 2258 1698 2262
rect 1750 2258 1754 2262
rect 1782 2258 1786 2262
rect 1838 2258 1842 2262
rect 1862 2258 1866 2262
rect 1894 2258 1898 2262
rect 1926 2258 1930 2262
rect 1942 2258 1946 2262
rect 1966 2258 1970 2262
rect 1974 2258 1978 2262
rect 2006 2258 2010 2262
rect 2022 2258 2026 2262
rect 2054 2258 2058 2262
rect 2078 2258 2082 2262
rect 2102 2258 2106 2262
rect 2126 2258 2130 2262
rect 2133 2258 2137 2262
rect 2270 2258 2274 2262
rect 2310 2258 2314 2262
rect 2334 2258 2338 2262
rect 2350 2258 2354 2262
rect 2366 2258 2370 2262
rect 2390 2258 2394 2262
rect 2406 2258 2410 2262
rect 2422 2258 2426 2262
rect 2470 2258 2474 2262
rect 2566 2258 2570 2262
rect 2582 2258 2586 2262
rect 2598 2258 2602 2262
rect 2606 2258 2610 2262
rect 2630 2258 2634 2262
rect 2798 2258 2802 2262
rect 2990 2258 2994 2262
rect 3134 2258 3138 2262
rect 3182 2258 3186 2262
rect 3206 2258 3210 2262
rect 3222 2258 3226 2262
rect 3238 2258 3242 2262
rect 3262 2258 3266 2262
rect 3286 2258 3290 2262
rect 3294 2258 3298 2262
rect 3326 2258 3330 2262
rect 3350 2258 3354 2262
rect 3358 2258 3362 2262
rect 3382 2258 3386 2262
rect 3398 2258 3402 2262
rect 3446 2258 3450 2262
rect 3478 2258 3482 2262
rect 3526 2258 3530 2262
rect 3558 2258 3562 2262
rect 3622 2258 3626 2262
rect 3638 2258 3642 2262
rect 3662 2258 3666 2262
rect 3670 2258 3674 2262
rect 3710 2258 3714 2262
rect 3742 2258 3746 2262
rect 3758 2258 3762 2262
rect 3766 2258 3770 2262
rect 3790 2258 3794 2262
rect 3846 2258 3850 2262
rect 3894 2258 3898 2262
rect 3934 2258 3938 2262
rect 3950 2258 3954 2262
rect 4006 2258 4010 2262
rect 4014 2258 4018 2262
rect 4030 2258 4034 2262
rect 4046 2258 4050 2262
rect 4086 2258 4090 2262
rect 4166 2258 4170 2262
rect 4198 2258 4202 2262
rect 4246 2258 4250 2262
rect 4270 2258 4274 2262
rect 4294 2258 4298 2262
rect 4318 2258 4322 2262
rect 4374 2258 4378 2262
rect 462 2248 466 2252
rect 486 2250 490 2254
rect 670 2248 674 2252
rect 702 2248 706 2252
rect 750 2248 754 2252
rect 782 2248 786 2252
rect 790 2248 794 2252
rect 814 2248 818 2252
rect 846 2248 850 2252
rect 878 2248 882 2252
rect 934 2248 938 2252
rect 1006 2248 1010 2252
rect 1094 2248 1098 2252
rect 1158 2250 1162 2254
rect 1318 2248 1322 2252
rect 1342 2248 1346 2252
rect 1390 2248 1394 2252
rect 1758 2248 1762 2252
rect 1870 2248 1874 2252
rect 1910 2248 1914 2252
rect 2022 2248 2026 2252
rect 2070 2248 2074 2252
rect 2262 2250 2266 2254
rect 2382 2248 2386 2252
rect 2486 2248 2490 2252
rect 2502 2248 2506 2252
rect 2550 2248 2554 2252
rect 2566 2248 2570 2252
rect 2782 2250 2786 2254
rect 2990 2248 2994 2252
rect 3166 2250 3170 2254
rect 3262 2248 3266 2252
rect 3318 2248 3322 2252
rect 3542 2248 3546 2252
rect 3558 2248 3562 2252
rect 3582 2248 3586 2252
rect 3646 2248 3650 2252
rect 3662 2248 3666 2252
rect 3726 2248 3730 2252
rect 3734 2248 3738 2252
rect 3822 2248 3826 2252
rect 3854 2248 3858 2252
rect 3878 2248 3882 2252
rect 3966 2248 3970 2252
rect 4062 2248 4066 2252
rect 4150 2248 4154 2252
rect 38 2238 42 2242
rect 798 2238 802 2242
rect 862 2238 866 2242
rect 1366 2238 1370 2242
rect 1678 2238 1682 2242
rect 1958 2238 1962 2242
rect 1974 2238 1978 2242
rect 3038 2238 3042 2242
rect 3526 2238 3530 2242
rect 3838 2238 3842 2242
rect 3902 2238 3906 2242
rect 3934 2238 3938 2242
rect 4126 2238 4130 2242
rect 54 2228 58 2232
rect 486 2227 490 2231
rect 1158 2227 1162 2231
rect 2262 2227 2266 2231
rect 2782 2227 2786 2231
rect 3166 2227 3170 2231
rect 3446 2228 3450 2232
rect 238 2218 242 2222
rect 270 2218 274 2222
rect 398 2218 402 2222
rect 614 2218 618 2222
rect 638 2218 642 2222
rect 966 2218 970 2222
rect 1062 2218 1066 2222
rect 1286 2218 1290 2222
rect 1390 2218 1394 2222
rect 1534 2218 1538 2222
rect 1766 2218 1770 2222
rect 1830 2218 1834 2222
rect 1846 2218 1850 2222
rect 2054 2218 2058 2222
rect 2086 2218 2090 2222
rect 2622 2218 2626 2222
rect 2654 2218 2658 2222
rect 2846 2218 2850 2222
rect 2990 2218 2994 2222
rect 3278 2218 3282 2222
rect 3846 2218 3850 2222
rect 3910 2218 3914 2222
rect 3950 2218 3954 2222
rect 4046 2218 4050 2222
rect 4350 2218 4354 2222
rect 394 2203 398 2207
rect 401 2203 405 2207
rect 1418 2203 1422 2207
rect 1425 2203 1429 2207
rect 2442 2203 2446 2207
rect 2449 2203 2453 2207
rect 3474 2203 3478 2207
rect 3481 2203 3485 2207
rect 54 2188 58 2192
rect 230 2188 234 2192
rect 366 2188 370 2192
rect 510 2188 514 2192
rect 678 2188 682 2192
rect 750 2188 754 2192
rect 774 2188 778 2192
rect 806 2188 810 2192
rect 870 2188 874 2192
rect 1014 2188 1018 2192
rect 1070 2188 1074 2192
rect 1150 2188 1154 2192
rect 1294 2188 1298 2192
rect 1462 2188 1466 2192
rect 1646 2188 1650 2192
rect 2206 2188 2210 2192
rect 2574 2188 2578 2192
rect 2726 2188 2730 2192
rect 2870 2188 2874 2192
rect 3302 2188 3306 2192
rect 3422 2188 3426 2192
rect 3590 2188 3594 2192
rect 3614 2188 3618 2192
rect 3694 2188 3698 2192
rect 3910 2188 3914 2192
rect 3958 2188 3962 2192
rect 3998 2188 4002 2192
rect 4030 2188 4034 2192
rect 4358 2188 4362 2192
rect 838 2178 842 2182
rect 6 2168 10 2172
rect 30 2168 34 2172
rect 718 2168 722 2172
rect 742 2168 746 2172
rect 814 2168 818 2172
rect 846 2168 850 2172
rect 862 2168 866 2172
rect 878 2168 882 2172
rect 950 2168 954 2172
rect 1806 2178 1810 2182
rect 2278 2178 2282 2182
rect 3126 2179 3130 2183
rect 3230 2178 3234 2182
rect 3406 2178 3410 2182
rect 4150 2178 4154 2182
rect 1366 2168 1370 2172
rect 1782 2168 1786 2172
rect 1814 2168 1818 2172
rect 2094 2168 2098 2172
rect 2998 2168 3002 2172
rect 4198 2168 4202 2172
rect 230 2158 234 2162
rect 254 2158 258 2162
rect 310 2158 314 2162
rect 366 2158 370 2162
rect 678 2158 682 2162
rect 758 2158 762 2162
rect 790 2158 794 2162
rect 798 2158 802 2162
rect 830 2158 834 2162
rect 862 2158 866 2162
rect 934 2158 938 2162
rect 966 2158 970 2162
rect 1118 2158 1122 2162
rect 1294 2158 1298 2162
rect 1350 2158 1354 2162
rect 1382 2158 1386 2162
rect 1422 2158 1426 2162
rect 1462 2158 1466 2162
rect 1686 2158 1690 2162
rect 1766 2158 1770 2162
rect 1798 2158 1802 2162
rect 1918 2158 1922 2162
rect 1982 2158 1986 2162
rect 2014 2158 2018 2162
rect 2046 2158 2050 2162
rect 2142 2158 2146 2162
rect 2198 2158 2202 2162
rect 2318 2158 2322 2162
rect 2350 2158 2354 2162
rect 2422 2158 2426 2162
rect 2566 2158 2570 2162
rect 2678 2158 2682 2162
rect 2870 2158 2874 2162
rect 2910 2158 2914 2162
rect 3126 2156 3130 2160
rect 3374 2158 3378 2162
rect 3726 2158 3730 2162
rect 3750 2158 3754 2162
rect 3774 2158 3778 2162
rect 3798 2158 3802 2162
rect 3886 2158 3890 2162
rect 4086 2158 4090 2162
rect 4134 2158 4138 2162
rect 4166 2158 4170 2162
rect 4214 2158 4218 2162
rect 4230 2158 4234 2162
rect 4270 2158 4274 2162
rect 22 2148 26 2152
rect 46 2148 50 2152
rect 70 2148 74 2152
rect 85 2148 89 2152
rect 222 2148 226 2152
rect 230 2148 234 2152
rect 262 2148 266 2152
rect 294 2148 298 2152
rect 310 2148 314 2152
rect 334 2148 338 2152
rect 374 2148 378 2152
rect 574 2148 578 2152
rect 702 2148 706 2152
rect 750 2148 754 2152
rect 774 2148 778 2152
rect 806 2148 810 2152
rect 838 2148 842 2152
rect 870 2148 874 2152
rect 918 2148 922 2152
rect 950 2148 954 2152
rect 998 2148 1002 2152
rect 1014 2148 1018 2152
rect 1030 2148 1034 2152
rect 1054 2148 1058 2152
rect 1070 2148 1074 2152
rect 1110 2148 1114 2152
rect 1118 2148 1122 2152
rect 1190 2148 1194 2152
rect 1246 2148 1250 2152
rect 1318 2148 1322 2152
rect 1358 2148 1362 2152
rect 1398 2148 1402 2152
rect 1510 2148 1514 2152
rect 1566 2148 1570 2152
rect 1622 2148 1626 2152
rect 1654 2148 1658 2152
rect 1662 2148 1666 2152
rect 1694 2148 1698 2152
rect 1702 2148 1706 2152
rect 1742 2148 1746 2152
rect 1758 2148 1762 2152
rect 1774 2148 1778 2152
rect 1806 2148 1810 2152
rect 1854 2148 1858 2152
rect 1862 2148 1866 2152
rect 1902 2148 1906 2152
rect 1950 2148 1954 2152
rect 1966 2148 1970 2152
rect 1982 2148 1986 2152
rect 1998 2148 2002 2152
rect 2022 2148 2026 2152
rect 2038 2148 2042 2152
rect 2062 2148 2066 2152
rect 2110 2148 2114 2152
rect 2126 2148 2130 2152
rect 2158 2148 2162 2152
rect 2174 2148 2178 2152
rect 2246 2148 2250 2152
rect 2302 2148 2306 2152
rect 2326 2148 2330 2152
rect 2358 2148 2362 2152
rect 2398 2148 2402 2152
rect 2438 2148 2442 2152
rect 2494 2148 2498 2152
rect 2558 2148 2562 2152
rect 2590 2148 2594 2152
rect 2598 2148 2602 2152
rect 2686 2148 2690 2152
rect 2854 2148 2858 2152
rect 2926 2148 2930 2152
rect 2958 2148 2962 2152
rect 3134 2148 3138 2152
rect 3190 2148 3194 2152
rect 3206 2148 3210 2152
rect 3238 2148 3242 2152
rect 3254 2148 3258 2152
rect 3270 2148 3274 2152
rect 3278 2148 3282 2152
rect 3310 2148 3314 2152
rect 3342 2148 3346 2152
rect 3358 2148 3362 2152
rect 3382 2148 3386 2152
rect 3422 2148 3426 2152
rect 3470 2148 3474 2152
rect 3494 2148 3498 2152
rect 3502 2148 3506 2152
rect 3526 2148 3530 2152
rect 3566 2148 3570 2152
rect 3574 2148 3578 2152
rect 3630 2148 3634 2152
rect 3750 2148 3754 2152
rect 3806 2148 3810 2152
rect 3838 2148 3842 2152
rect 3894 2148 3898 2152
rect 3926 2148 3930 2152
rect 4014 2148 4018 2152
rect 4046 2148 4050 2152
rect 182 2138 186 2142
rect 286 2138 290 2142
rect 318 2138 322 2142
rect 414 2138 418 2142
rect 533 2138 537 2142
rect 630 2138 634 2142
rect 766 2138 770 2142
rect 910 2138 914 2142
rect 926 2138 930 2142
rect 942 2138 946 2142
rect 1006 2138 1010 2142
rect 1038 2138 1042 2142
rect 1046 2138 1050 2142
rect 1078 2138 1082 2142
rect 1086 2138 1090 2142
rect 1142 2138 1146 2142
rect 1246 2138 1250 2142
rect 1318 2138 1322 2142
rect 1334 2138 1338 2142
rect 1414 2138 1418 2142
rect 1510 2138 1514 2142
rect 1630 2138 1634 2142
rect 1646 2138 1650 2142
rect 1662 2138 1666 2142
rect 1686 2138 1690 2142
rect 1710 2138 1714 2142
rect 1718 2138 1722 2142
rect 1726 2138 1730 2142
rect 1758 2138 1762 2142
rect 1894 2138 1898 2142
rect 1942 2138 1946 2142
rect 1958 2138 1962 2142
rect 1982 2138 1986 2142
rect 2006 2138 2010 2142
rect 2038 2138 2042 2142
rect 2054 2138 2058 2142
rect 2070 2138 2074 2142
rect 2078 2138 2082 2142
rect 2094 2138 2098 2142
rect 2118 2138 2122 2142
rect 2166 2138 2170 2142
rect 2174 2138 2178 2142
rect 2254 2138 2258 2142
rect 2294 2138 2298 2142
rect 2326 2138 2330 2142
rect 2382 2138 2386 2142
rect 2390 2138 2394 2142
rect 2430 2138 2434 2142
rect 2446 2138 2450 2142
rect 2454 2138 2458 2142
rect 2502 2138 2506 2142
rect 2582 2138 2586 2142
rect 2630 2138 2634 2142
rect 2638 2138 2642 2142
rect 2654 2138 2658 2142
rect 2694 2138 2698 2142
rect 2822 2138 2826 2142
rect 2894 2138 2898 2142
rect 2902 2138 2906 2142
rect 2934 2138 2938 2142
rect 2982 2138 2986 2142
rect 3094 2138 3098 2142
rect 3166 2138 3170 2142
rect 3182 2138 3186 2142
rect 3214 2138 3218 2142
rect 3246 2138 3250 2142
rect 3262 2138 3266 2142
rect 3286 2138 3290 2142
rect 3318 2138 3322 2142
rect 3334 2138 3338 2142
rect 3350 2138 3354 2142
rect 3366 2138 3370 2142
rect 3390 2138 3394 2142
rect 3414 2138 3418 2142
rect 3462 2138 3466 2142
rect 3534 2138 3538 2142
rect 3638 2138 3642 2142
rect 3710 2138 3714 2142
rect 3734 2138 3738 2142
rect 4102 2148 4106 2152
rect 4150 2148 4154 2152
rect 4190 2148 4194 2152
rect 4230 2148 4234 2152
rect 4254 2148 4258 2152
rect 3758 2138 3762 2142
rect 3774 2138 3778 2142
rect 3782 2138 3786 2142
rect 3830 2138 3834 2142
rect 3870 2138 3874 2142
rect 3886 2138 3890 2142
rect 3918 2138 3922 2142
rect 3966 2138 3970 2142
rect 4054 2138 4058 2142
rect 4062 2138 4066 2142
rect 4110 2138 4114 2142
rect 4118 2138 4122 2142
rect 4142 2138 4146 2142
rect 4238 2138 4242 2142
rect 4246 2138 4250 2142
rect 4278 2138 4282 2142
rect 4326 2138 4330 2142
rect 4382 2138 4386 2142
rect 166 2128 170 2132
rect 430 2128 434 2132
rect 526 2128 530 2132
rect 614 2128 618 2132
rect 1230 2128 1234 2132
rect 1390 2128 1394 2132
rect 1526 2128 1530 2132
rect 1614 2128 1618 2132
rect 1742 2128 1746 2132
rect 2086 2128 2090 2132
rect 2214 2128 2218 2132
rect 2470 2128 2474 2132
rect 2502 2128 2506 2132
rect 2534 2128 2538 2132
rect 2558 2128 2562 2132
rect 2710 2128 2714 2132
rect 2806 2128 2810 2132
rect 3078 2128 3082 2132
rect 3166 2128 3170 2132
rect 3406 2128 3410 2132
rect 3446 2128 3450 2132
rect 3830 2128 3834 2132
rect 3862 2128 3866 2132
rect 4070 2128 4074 2132
rect 4078 2128 4082 2132
rect 4174 2128 4178 2132
rect 982 2118 986 2122
rect 1782 2118 1786 2122
rect 1838 2118 1842 2122
rect 1878 2118 1882 2122
rect 1918 2118 1922 2122
rect 2198 2118 2202 2122
rect 2230 2118 2234 2122
rect 2318 2118 2322 2122
rect 2350 2118 2354 2122
rect 2414 2118 2418 2122
rect 2646 2118 2650 2122
rect 2678 2118 2682 2122
rect 2702 2118 2706 2122
rect 2910 2118 2914 2122
rect 3198 2118 3202 2122
rect 3326 2118 3330 2122
rect 3550 2118 3554 2122
rect 3614 2118 3618 2122
rect 3726 2118 3730 2122
rect 3822 2118 3826 2122
rect 3854 2118 3858 2122
rect 3942 2118 3946 2122
rect 4086 2118 4090 2122
rect 4134 2118 4138 2122
rect 4270 2118 4274 2122
rect 4294 2118 4298 2122
rect 898 2103 902 2107
rect 905 2103 909 2107
rect 1930 2103 1934 2107
rect 1937 2103 1941 2107
rect 2954 2103 2958 2107
rect 2961 2103 2965 2107
rect 3978 2103 3982 2107
rect 3985 2103 3989 2107
rect 518 2088 522 2092
rect 550 2088 554 2092
rect 678 2088 682 2092
rect 686 2088 690 2092
rect 766 2088 770 2092
rect 838 2088 842 2092
rect 886 2088 890 2092
rect 918 2088 922 2092
rect 974 2088 978 2092
rect 1070 2088 1074 2092
rect 1446 2088 1450 2092
rect 1486 2088 1490 2092
rect 1598 2088 1602 2092
rect 2078 2088 2082 2092
rect 2182 2088 2186 2092
rect 2382 2088 2386 2092
rect 2406 2088 2410 2092
rect 2526 2088 2530 2092
rect 2838 2088 2842 2092
rect 3262 2088 3266 2092
rect 3294 2088 3298 2092
rect 3462 2088 3466 2092
rect 3486 2088 3490 2092
rect 3566 2088 3570 2092
rect 3582 2088 3586 2092
rect 3606 2088 3610 2092
rect 3870 2088 3874 2092
rect 4070 2088 4074 2092
rect 4150 2088 4154 2092
rect 4278 2088 4282 2092
rect 4382 2088 4386 2092
rect 166 2078 170 2082
rect 334 2078 338 2082
rect 646 2078 650 2082
rect 726 2078 730 2082
rect 1286 2078 1290 2082
rect 1382 2078 1386 2082
rect 1710 2078 1714 2082
rect 1806 2078 1810 2082
rect 1966 2078 1970 2082
rect 2006 2078 2010 2082
rect 2046 2078 2050 2082
rect 2110 2078 2114 2082
rect 2126 2078 2130 2082
rect 2286 2078 2290 2082
rect 2390 2078 2394 2082
rect 2622 2078 2626 2082
rect 2870 2078 2874 2082
rect 3086 2078 3090 2082
rect 3230 2078 3234 2082
rect 3358 2078 3362 2082
rect 3470 2078 3474 2082
rect 3526 2078 3530 2082
rect 3734 2078 3738 2082
rect 3830 2078 3834 2082
rect 3918 2078 3922 2082
rect 3934 2078 3938 2082
rect 4078 2078 4082 2082
rect 4190 2078 4194 2082
rect 4246 2078 4250 2082
rect 4390 2078 4394 2082
rect 54 2068 58 2072
rect 85 2068 89 2072
rect 182 2068 186 2072
rect 318 2068 322 2072
rect 446 2068 450 2072
rect 462 2068 466 2072
rect 494 2068 498 2072
rect 534 2068 538 2072
rect 606 2068 610 2072
rect 614 2068 618 2072
rect 654 2068 658 2072
rect 710 2068 714 2072
rect 718 2068 722 2072
rect 790 2068 794 2072
rect 862 2068 866 2072
rect 942 2068 946 2072
rect 998 2068 1002 2072
rect 1006 2068 1010 2072
rect 1038 2068 1042 2072
rect 1046 2068 1050 2072
rect 1102 2068 1106 2072
rect 1134 2068 1138 2072
rect 1182 2068 1186 2072
rect 1198 2068 1202 2072
rect 1270 2068 1274 2072
rect 1406 2068 1410 2072
rect 1462 2068 1466 2072
rect 1494 2068 1498 2072
rect 1590 2068 1594 2072
rect 1606 2068 1610 2072
rect 1622 2068 1626 2072
rect 1726 2068 1730 2072
rect 1838 2068 1842 2072
rect 1846 2068 1850 2072
rect 1878 2068 1882 2072
rect 1918 2068 1922 2072
rect 1958 2068 1962 2072
rect 1982 2068 1986 2072
rect 2014 2068 2018 2072
rect 2110 2068 2114 2072
rect 2158 2068 2162 2072
rect 2302 2068 2306 2072
rect 2398 2068 2402 2072
rect 2430 2068 2434 2072
rect 2454 2068 2458 2072
rect 2470 2068 2474 2072
rect 2502 2068 2506 2072
rect 2638 2068 2642 2072
rect 2710 2068 2714 2072
rect 2734 2068 2738 2072
rect 2742 2068 2746 2072
rect 2774 2068 2778 2072
rect 2798 2068 2802 2072
rect 2830 2068 2834 2072
rect 2862 2068 2866 2072
rect 2894 2068 2898 2072
rect 2902 2068 2906 2072
rect 2934 2068 2938 2072
rect 2950 2068 2954 2072
rect 3102 2068 3106 2072
rect 3182 2068 3186 2072
rect 3198 2068 3202 2072
rect 3206 2068 3210 2072
rect 3238 2068 3242 2072
rect 3270 2068 3274 2072
rect 3286 2068 3290 2072
rect 3334 2068 3338 2072
rect 3422 2068 3426 2072
rect 3438 2068 3442 2072
rect 3454 2068 3458 2072
rect 3518 2068 3522 2072
rect 3542 2068 3546 2072
rect 3574 2068 3578 2072
rect 3598 2068 3602 2072
rect 3630 2068 3634 2072
rect 3646 2068 3650 2072
rect 3686 2068 3690 2072
rect 3718 2068 3722 2072
rect 3766 2068 3770 2072
rect 3782 2068 3786 2072
rect 3798 2068 3802 2072
rect 3894 2068 3898 2072
rect 4006 2068 4010 2072
rect 4030 2068 4034 2072
rect 4118 2068 4122 2072
rect 4174 2068 4178 2072
rect 4206 2068 4210 2072
rect 4238 2068 4242 2072
rect 4326 2068 4330 2072
rect 4358 2068 4362 2072
rect 46 2058 50 2062
rect 62 2058 66 2062
rect 230 2058 234 2062
rect 270 2058 274 2062
rect 374 2058 378 2062
rect 470 2058 474 2062
rect 486 2058 490 2062
rect 502 2058 506 2062
rect 518 2058 522 2062
rect 630 2058 634 2062
rect 662 2058 666 2062
rect 702 2058 706 2062
rect 750 2058 754 2062
rect 782 2058 786 2062
rect 806 2058 810 2062
rect 854 2058 858 2062
rect 870 2058 874 2062
rect 934 2058 938 2062
rect 942 2058 946 2062
rect 958 2058 962 2062
rect 990 2058 994 2062
rect 1006 2058 1010 2062
rect 1030 2058 1034 2062
rect 1054 2058 1058 2062
rect 1078 2058 1082 2062
rect 1126 2058 1130 2062
rect 1150 2058 1154 2062
rect 1198 2058 1202 2062
rect 1222 2058 1226 2062
rect 1398 2058 1402 2062
rect 1406 2058 1410 2062
rect 1470 2058 1474 2062
rect 1566 2058 1570 2062
rect 1766 2058 1770 2062
rect 1806 2058 1810 2062
rect 1830 2058 1834 2062
rect 1854 2058 1858 2062
rect 1870 2058 1874 2062
rect 1886 2058 1890 2062
rect 1902 2058 1906 2062
rect 1950 2058 1954 2062
rect 1990 2058 1994 2062
rect 2022 2058 2026 2062
rect 2038 2058 2042 2062
rect 2062 2058 2066 2062
rect 2078 2058 2082 2062
rect 2102 2058 2106 2062
rect 2110 2058 2114 2062
rect 2126 2058 2130 2062
rect 2150 2058 2154 2062
rect 2166 2058 2170 2062
rect 2334 2058 2338 2062
rect 2374 2058 2378 2062
rect 2422 2058 2426 2062
rect 2438 2058 2442 2062
rect 2478 2058 2482 2062
rect 2582 2058 2586 2062
rect 2726 2058 2730 2062
rect 2742 2058 2746 2062
rect 2798 2058 2802 2062
rect 2838 2058 2842 2062
rect 2854 2058 2858 2062
rect 2886 2058 2890 2062
rect 2910 2058 2914 2062
rect 2926 2058 2930 2062
rect 2990 2058 2994 2062
rect 3046 2058 3050 2062
rect 3134 2058 3138 2062
rect 3190 2058 3194 2062
rect 3214 2058 3218 2062
rect 3246 2058 3250 2062
rect 3262 2058 3266 2062
rect 3278 2058 3282 2062
rect 3326 2058 3330 2062
rect 3342 2058 3346 2062
rect 3366 2058 3370 2062
rect 3374 2058 3378 2062
rect 3398 2058 3402 2062
rect 3406 2058 3410 2062
rect 3430 2058 3434 2062
rect 3446 2058 3450 2062
rect 3510 2058 3514 2062
rect 3550 2058 3554 2062
rect 3622 2058 3626 2062
rect 3646 2058 3650 2062
rect 3654 2058 3658 2062
rect 3678 2058 3682 2062
rect 3710 2058 3714 2062
rect 3758 2058 3762 2062
rect 3774 2058 3778 2062
rect 3806 2058 3810 2062
rect 3814 2058 3818 2062
rect 3846 2058 3850 2062
rect 3854 2058 3858 2062
rect 3878 2058 3882 2062
rect 3918 2058 3922 2062
rect 4054 2058 4058 2062
rect 4102 2058 4106 2062
rect 4126 2058 4130 2062
rect 4166 2058 4170 2062
rect 4206 2058 4210 2062
rect 4270 2058 4274 2062
rect 4302 2058 4306 2062
rect 4326 2058 4330 2062
rect 4350 2058 4354 2062
rect 30 2048 34 2052
rect 214 2050 218 2054
rect 286 2050 290 2054
rect 486 2048 490 2052
rect 518 2048 522 2052
rect 622 2048 626 2052
rect 678 2048 682 2052
rect 686 2048 690 2052
rect 734 2048 738 2052
rect 742 2048 746 2052
rect 766 2048 770 2052
rect 798 2048 802 2052
rect 886 2048 890 2052
rect 966 2048 970 2052
rect 974 2048 978 2052
rect 1070 2048 1074 2052
rect 1110 2048 1114 2052
rect 1142 2048 1146 2052
rect 1238 2050 1242 2054
rect 1366 2048 1370 2052
rect 1382 2048 1386 2052
rect 1486 2048 1490 2052
rect 1774 2048 1778 2052
rect 1814 2048 1818 2052
rect 1870 2048 1874 2052
rect 1934 2048 1938 2052
rect 2038 2048 2042 2052
rect 2134 2048 2138 2052
rect 2350 2048 2354 2052
rect 2494 2048 2498 2052
rect 2526 2048 2530 2052
rect 2670 2050 2674 2054
rect 2710 2048 2714 2052
rect 2750 2048 2754 2052
rect 2766 2048 2770 2052
rect 2782 2048 2786 2052
rect 2790 2048 2794 2052
rect 2806 2048 2810 2052
rect 2822 2048 2826 2052
rect 2926 2048 2930 2052
rect 3150 2048 3154 2052
rect 3174 2048 3178 2052
rect 3310 2048 3314 2052
rect 3414 2048 3418 2052
rect 3494 2048 3498 2052
rect 3558 2048 3562 2052
rect 3582 2048 3586 2052
rect 3606 2048 3610 2052
rect 3702 2048 3706 2052
rect 3758 2048 3762 2052
rect 3910 2048 3914 2052
rect 4046 2048 4050 2052
rect 4110 2048 4114 2052
rect 4142 2048 4146 2052
rect 4150 2048 4154 2052
rect 4262 2048 4266 2052
rect 4294 2048 4298 2052
rect 4334 2048 4338 2052
rect 6 2038 10 2042
rect 814 2038 818 2042
rect 1126 2038 1130 2042
rect 1158 2038 1162 2042
rect 1990 2038 1994 2042
rect 4094 2038 4098 2042
rect 4278 2038 4282 2042
rect 4310 2038 4314 2042
rect 286 2027 290 2031
rect 742 2028 746 2032
rect 1238 2027 1242 2031
rect 2542 2028 2546 2032
rect 2670 2027 2674 2031
rect 3526 2028 3530 2032
rect 4302 2028 4306 2032
rect 70 2018 74 2022
rect 214 2018 218 2022
rect 630 2018 634 2022
rect 806 2018 810 2022
rect 838 2018 842 2022
rect 1030 2018 1034 2022
rect 1550 2018 1554 2022
rect 1598 2018 1602 2022
rect 1630 2018 1634 2022
rect 1774 2018 1778 2022
rect 1798 2018 1802 2022
rect 1886 2018 1890 2022
rect 1950 2018 1954 2022
rect 2206 2018 2210 2022
rect 2350 2018 2354 2022
rect 2942 2018 2946 2022
rect 2974 2018 2978 2022
rect 3006 2018 3010 2022
rect 3150 2018 3154 2022
rect 3782 2018 3786 2022
rect 3918 2018 3922 2022
rect 3950 2018 3954 2022
rect 4102 2018 4106 2022
rect 4126 2018 4130 2022
rect 4254 2018 4258 2022
rect 4382 2018 4386 2022
rect 394 2003 398 2007
rect 401 2003 405 2007
rect 1418 2003 1422 2007
rect 1425 2003 1429 2007
rect 2442 2003 2446 2007
rect 2449 2003 2453 2007
rect 3474 2003 3478 2007
rect 3481 2003 3485 2007
rect 6 1988 10 1992
rect 30 1988 34 1992
rect 142 1988 146 1992
rect 398 1988 402 1992
rect 622 1988 626 1992
rect 694 1988 698 1992
rect 766 1988 770 1992
rect 830 1988 834 1992
rect 1022 1988 1026 1992
rect 1062 1988 1066 1992
rect 1174 1988 1178 1992
rect 1390 1988 1394 1992
rect 1486 1988 1490 1992
rect 1750 1988 1754 1992
rect 1830 1988 1834 1992
rect 1862 1988 1866 1992
rect 1966 1988 1970 1992
rect 2054 1988 2058 1992
rect 2230 1988 2234 1992
rect 2430 1988 2434 1992
rect 2614 1988 2618 1992
rect 2646 1988 2650 1992
rect 2670 1988 2674 1992
rect 2814 1988 2818 1992
rect 2846 1988 2850 1992
rect 2990 1988 2994 1992
rect 3294 1988 3298 1992
rect 3326 1988 3330 1992
rect 3630 1988 3634 1992
rect 3662 1988 3666 1992
rect 3686 1988 3690 1992
rect 3710 1988 3714 1992
rect 3910 1988 3914 1992
rect 4118 1988 4122 1992
rect 4230 1988 4234 1992
rect 4278 1988 4282 1992
rect 118 1978 122 1982
rect 574 1979 578 1983
rect 734 1978 738 1982
rect 862 1978 866 1982
rect 638 1968 642 1972
rect 702 1968 706 1972
rect 742 1968 746 1972
rect 774 1968 778 1972
rect 838 1968 842 1972
rect 926 1968 930 1972
rect 966 1968 970 1972
rect 1030 1968 1034 1972
rect 1054 1968 1058 1972
rect 1158 1968 1162 1972
rect 1262 1978 1266 1982
rect 1542 1979 1546 1983
rect 3278 1978 3282 1982
rect 3766 1978 3770 1982
rect 4150 1978 4154 1982
rect 1246 1968 1250 1972
rect 1302 1968 1306 1972
rect 1342 1968 1346 1972
rect 1494 1968 1498 1972
rect 2582 1968 2586 1972
rect 4142 1968 4146 1972
rect 4214 1968 4218 1972
rect 4238 1968 4242 1972
rect 4270 1968 4274 1972
rect 62 1958 66 1962
rect 78 1958 82 1962
rect 94 1958 98 1962
rect 110 1958 114 1962
rect 174 1958 178 1962
rect 190 1958 194 1962
rect 222 1958 226 1962
rect 238 1958 242 1962
rect 398 1958 402 1962
rect 574 1956 578 1960
rect 654 1958 658 1962
rect 686 1958 690 1962
rect 726 1958 730 1962
rect 758 1958 762 1962
rect 790 1958 794 1962
rect 822 1958 826 1962
rect 950 1958 954 1962
rect 982 1958 986 1962
rect 1014 1958 1018 1962
rect 1070 1958 1074 1962
rect 1166 1958 1170 1962
rect 1230 1958 1234 1962
rect 1278 1958 1282 1962
rect 1318 1958 1322 1962
rect 1478 1958 1482 1962
rect 22 1948 26 1952
rect 46 1948 50 1952
rect 62 1948 66 1952
rect 94 1948 98 1952
rect 134 1948 138 1952
rect 158 1948 162 1952
rect 174 1948 178 1952
rect 206 1948 210 1952
rect 230 1948 234 1952
rect 398 1948 402 1952
rect 590 1948 594 1952
rect 614 1948 618 1952
rect 638 1948 642 1952
rect 662 1948 666 1952
rect 686 1948 690 1952
rect 710 1948 714 1952
rect 734 1948 738 1952
rect 766 1948 770 1952
rect 814 1948 818 1952
rect 830 1948 834 1952
rect 878 1948 882 1952
rect 926 1948 930 1952
rect 958 1948 962 1952
rect 982 1948 986 1952
rect 998 1948 1002 1952
rect 1022 1948 1026 1952
rect 1062 1948 1066 1952
rect 1086 1948 1090 1952
rect 1102 1948 1106 1952
rect 1134 1948 1138 1952
rect 1174 1948 1178 1952
rect 1206 1948 1210 1952
rect 1238 1948 1242 1952
rect 1542 1956 1546 1960
rect 1718 1958 1722 1962
rect 1758 1958 1762 1962
rect 1942 1958 1946 1962
rect 1982 1958 1986 1962
rect 2014 1958 2018 1962
rect 2230 1958 2234 1962
rect 2430 1958 2434 1962
rect 2510 1958 2514 1962
rect 2542 1958 2546 1962
rect 2638 1958 2642 1962
rect 2814 1958 2818 1962
rect 2990 1958 2994 1962
rect 3054 1958 3058 1962
rect 3086 1958 3090 1962
rect 3102 1958 3106 1962
rect 3134 1958 3138 1962
rect 3198 1958 3202 1962
rect 3510 1958 3514 1962
rect 3550 1958 3554 1962
rect 3606 1958 3610 1962
rect 3910 1958 3914 1962
rect 3958 1958 3962 1962
rect 4014 1958 4018 1962
rect 4158 1958 4162 1962
rect 4198 1958 4202 1962
rect 4254 1958 4258 1962
rect 4286 1958 4290 1962
rect 4334 1958 4338 1962
rect 1302 1948 1306 1952
rect 1358 1948 1362 1952
rect 1382 1948 1386 1952
rect 1430 1948 1434 1952
rect 1438 1948 1442 1952
rect 1470 1948 1474 1952
rect 1486 1948 1490 1952
rect 1526 1948 1530 1952
rect 1678 1948 1682 1952
rect 1774 1948 1778 1952
rect 1782 1948 1786 1952
rect 1790 1948 1794 1952
rect 1846 1948 1850 1952
rect 1878 1948 1882 1952
rect 1934 1948 1938 1952
rect 2006 1948 2010 1952
rect 2038 1948 2042 1952
rect 2070 1948 2074 1952
rect 2126 1948 2130 1952
rect 2230 1948 2234 1952
rect 2270 1948 2274 1952
rect 2326 1948 2330 1952
rect 2430 1948 2434 1952
rect 2478 1948 2482 1952
rect 2494 1948 2498 1952
rect 2510 1948 2514 1952
rect 2558 1948 2562 1952
rect 2590 1948 2594 1952
rect 2598 1948 2602 1952
rect 2622 1948 2626 1952
rect 2814 1948 2818 1952
rect 54 1938 58 1942
rect 86 1938 90 1942
rect 166 1938 170 1942
rect 198 1938 202 1942
rect 214 1938 218 1942
rect 253 1938 257 1942
rect 350 1938 354 1942
rect 445 1938 449 1942
rect 542 1938 546 1942
rect 630 1938 634 1942
rect 662 1938 666 1942
rect 814 1938 818 1942
rect 886 1938 890 1942
rect 918 1938 922 1942
rect 2990 1948 2994 1952
rect 3014 1948 3018 1952
rect 3070 1948 3074 1952
rect 3102 1948 3106 1952
rect 3118 1948 3122 1952
rect 3134 1948 3138 1952
rect 3150 1948 3154 1952
rect 3190 1948 3194 1952
rect 3206 1948 3210 1952
rect 3214 1948 3218 1952
rect 3230 1948 3234 1952
rect 3254 1948 3258 1952
rect 3310 1948 3314 1952
rect 3342 1948 3346 1952
rect 3390 1948 3394 1952
rect 3406 1948 3410 1952
rect 3422 1948 3426 1952
rect 3430 1948 3434 1952
rect 3510 1948 3514 1952
rect 3518 1948 3522 1952
rect 3526 1948 3530 1952
rect 3550 1948 3554 1952
rect 3598 1948 3602 1952
rect 3630 1948 3634 1952
rect 3646 1948 3650 1952
rect 3694 1948 3698 1952
rect 3718 1948 3722 1952
rect 3726 1948 3730 1952
rect 3902 1948 3906 1952
rect 3950 1948 3954 1952
rect 4070 1948 4074 1952
rect 4094 1948 4098 1952
rect 4102 1948 4106 1952
rect 4150 1948 4154 1952
rect 4166 1948 4170 1952
rect 4198 1948 4202 1952
rect 4214 1948 4218 1952
rect 4246 1948 4250 1952
rect 4278 1948 4282 1952
rect 4366 1948 4370 1952
rect 1006 1938 1010 1942
rect 1078 1938 1082 1942
rect 1110 1938 1114 1942
rect 1142 1938 1146 1942
rect 1158 1938 1162 1942
rect 1198 1938 1202 1942
rect 1270 1938 1274 1942
rect 1326 1938 1330 1942
rect 1350 1938 1354 1942
rect 1382 1938 1386 1942
rect 1406 1938 1410 1942
rect 1446 1938 1450 1942
rect 1462 1938 1466 1942
rect 1574 1938 1578 1942
rect 1694 1938 1698 1942
rect 1718 1938 1722 1942
rect 1734 1938 1738 1942
rect 1742 1938 1746 1942
rect 1758 1938 1762 1942
rect 1798 1938 1802 1942
rect 1806 1938 1810 1942
rect 1910 1938 1914 1942
rect 1998 1938 2002 1942
rect 2014 1938 2018 1942
rect 2046 1938 2050 1942
rect 2182 1938 2186 1942
rect 2382 1938 2386 1942
rect 2462 1938 2466 1942
rect 2486 1938 2490 1942
rect 2502 1938 2506 1942
rect 2534 1938 2538 1942
rect 2566 1938 2570 1942
rect 2654 1938 2658 1942
rect 2766 1938 2770 1942
rect 2886 1938 2890 1942
rect 2942 1938 2946 1942
rect 3030 1938 3034 1942
rect 3062 1938 3066 1942
rect 3094 1938 3098 1942
rect 3126 1938 3130 1942
rect 3158 1938 3162 1942
rect 3182 1938 3186 1942
rect 3222 1938 3226 1942
rect 3262 1938 3266 1942
rect 3350 1938 3354 1942
rect 3398 1938 3402 1942
rect 3414 1938 3418 1942
rect 3438 1938 3442 1942
rect 3454 1938 3458 1942
rect 3534 1938 3538 1942
rect 3542 1938 3546 1942
rect 3590 1938 3594 1942
rect 3622 1938 3626 1942
rect 3678 1938 3682 1942
rect 3862 1938 3866 1942
rect 3974 1938 3978 1942
rect 4014 1938 4018 1942
rect 4174 1938 4178 1942
rect 4222 1938 4226 1942
rect 4294 1938 4298 1942
rect 4318 1938 4322 1942
rect 4358 1938 4362 1942
rect 334 1928 338 1932
rect 526 1928 530 1932
rect 1086 1928 1090 1932
rect 1118 1928 1122 1932
rect 1278 1928 1282 1932
rect 1358 1928 1362 1932
rect 1390 1928 1394 1932
rect 1590 1928 1594 1932
rect 1710 1928 1714 1932
rect 1958 1928 1962 1932
rect 1974 1928 1978 1932
rect 2078 1928 2082 1932
rect 2166 1928 2170 1932
rect 2254 1928 2258 1932
rect 2278 1928 2282 1932
rect 2366 1928 2370 1932
rect 2574 1928 2578 1932
rect 2750 1928 2754 1932
rect 2926 1928 2930 1932
rect 3054 1928 3058 1932
rect 3086 1928 3090 1932
rect 3166 1928 3170 1932
rect 3246 1928 3250 1932
rect 3278 1928 3282 1932
rect 3574 1928 3578 1932
rect 3654 1928 3658 1932
rect 3678 1928 3682 1932
rect 3702 1928 3706 1932
rect 3846 1928 3850 1932
rect 3934 1928 3938 1932
rect 4022 1928 4026 1932
rect 4038 1928 4042 1932
rect 4070 1928 4074 1932
rect 4190 1928 4194 1932
rect 4294 1928 4298 1932
rect 4342 1928 4346 1932
rect 790 1918 794 1922
rect 1222 1918 1226 1922
rect 1334 1918 1338 1922
rect 1454 1918 1458 1922
rect 1670 1918 1674 1922
rect 1726 1918 1730 1922
rect 1814 1918 1818 1922
rect 1894 1918 1898 1922
rect 1942 1918 1946 1922
rect 1990 1918 1994 1922
rect 2054 1918 2058 1922
rect 2262 1918 2266 1922
rect 3174 1918 3178 1922
rect 3358 1918 3362 1922
rect 3446 1918 3450 1922
rect 3742 1918 3746 1922
rect 3942 1918 3946 1922
rect 3958 1918 3962 1922
rect 4006 1918 4010 1922
rect 4046 1918 4050 1922
rect 4062 1918 4066 1922
rect 4086 1918 4090 1922
rect 4334 1918 4338 1922
rect 4350 1918 4354 1922
rect 898 1903 902 1907
rect 905 1903 909 1907
rect 1930 1903 1934 1907
rect 1937 1903 1941 1907
rect 2954 1903 2958 1907
rect 2961 1903 2965 1907
rect 3978 1903 3982 1907
rect 3985 1903 3989 1907
rect 286 1888 290 1892
rect 630 1888 634 1892
rect 742 1888 746 1892
rect 958 1888 962 1892
rect 974 1888 978 1892
rect 1062 1888 1066 1892
rect 1190 1888 1194 1892
rect 1310 1888 1314 1892
rect 1446 1888 1450 1892
rect 1478 1888 1482 1892
rect 1534 1888 1538 1892
rect 1606 1888 1610 1892
rect 1638 1888 1642 1892
rect 1774 1888 1778 1892
rect 1998 1888 2002 1892
rect 2022 1888 2026 1892
rect 2230 1888 2234 1892
rect 2374 1888 2378 1892
rect 2462 1888 2466 1892
rect 2710 1888 2714 1892
rect 2870 1888 2874 1892
rect 3062 1888 3066 1892
rect 3134 1888 3138 1892
rect 3174 1888 3178 1892
rect 3278 1888 3282 1892
rect 3534 1888 3538 1892
rect 3702 1888 3706 1892
rect 3726 1888 3730 1892
rect 4278 1888 4282 1892
rect 4302 1888 4306 1892
rect 174 1878 178 1882
rect 366 1878 370 1882
rect 550 1878 554 1882
rect 870 1878 874 1882
rect 1238 1878 1242 1882
rect 1510 1878 1514 1882
rect 1574 1878 1578 1882
rect 1646 1878 1650 1882
rect 1750 1878 1754 1882
rect 1766 1878 1770 1882
rect 1782 1878 1786 1882
rect 1870 1878 1874 1882
rect 2014 1878 2018 1882
rect 2222 1878 2226 1882
rect 2358 1878 2362 1882
rect 2390 1878 2394 1882
rect 2398 1878 2402 1882
rect 2590 1878 2594 1882
rect 2678 1878 2682 1882
rect 2742 1878 2746 1882
rect 3142 1878 3146 1882
rect 3414 1878 3418 1882
rect 3622 1878 3626 1882
rect 3710 1878 3714 1882
rect 3806 1878 3810 1882
rect 3878 1878 3882 1882
rect 3998 1878 4002 1882
rect 4046 1878 4050 1882
rect 4086 1878 4090 1882
rect 4102 1878 4106 1882
rect 4238 1878 4242 1882
rect 4310 1878 4314 1882
rect 4382 1878 4386 1882
rect 30 1868 34 1872
rect 54 1868 58 1872
rect 190 1868 194 1872
rect 262 1868 266 1872
rect 382 1868 386 1872
rect 534 1868 538 1872
rect 638 1868 642 1872
rect 734 1868 738 1872
rect 766 1868 770 1872
rect 774 1868 778 1872
rect 806 1868 810 1872
rect 822 1868 826 1872
rect 846 1868 850 1872
rect 878 1868 882 1872
rect 886 1868 890 1872
rect 902 1868 906 1872
rect 926 1868 930 1872
rect 966 1868 970 1872
rect 998 1868 1002 1872
rect 1006 1868 1010 1872
rect 1038 1868 1042 1872
rect 1094 1868 1098 1872
rect 1158 1868 1162 1872
rect 1166 1868 1170 1872
rect 1198 1868 1202 1872
rect 1214 1868 1218 1872
rect 1278 1868 1282 1872
rect 1294 1868 1298 1872
rect 1334 1868 1338 1872
rect 1342 1868 1346 1872
rect 1374 1868 1378 1872
rect 1470 1868 1474 1872
rect 1502 1868 1506 1872
rect 1550 1868 1554 1872
rect 1566 1868 1570 1872
rect 1614 1868 1618 1872
rect 1630 1868 1634 1872
rect 1654 1868 1658 1872
rect 1686 1868 1690 1872
rect 1710 1868 1714 1872
rect 1726 1868 1730 1872
rect 1742 1868 1746 1872
rect 1854 1868 1858 1872
rect 2014 1868 2018 1872
rect 2030 1868 2034 1872
rect 2054 1868 2058 1872
rect 2062 1868 2066 1872
rect 2094 1868 2098 1872
rect 2246 1868 2250 1872
rect 2254 1866 2258 1870
rect 22 1858 26 1862
rect 54 1858 58 1862
rect 62 1858 66 1862
rect 78 1858 82 1862
rect 190 1858 194 1862
rect 246 1858 250 1862
rect 382 1858 386 1862
rect 430 1858 434 1862
rect 78 1848 82 1852
rect 94 1848 98 1852
rect 238 1848 242 1852
rect 278 1848 282 1852
rect 414 1850 418 1854
rect 590 1858 594 1862
rect 654 1858 658 1862
rect 662 1858 666 1862
rect 694 1858 698 1862
rect 710 1858 714 1862
rect 726 1858 730 1862
rect 758 1858 762 1862
rect 782 1858 786 1862
rect 814 1858 818 1862
rect 830 1858 834 1862
rect 854 1858 858 1862
rect 870 1858 874 1862
rect 894 1858 898 1862
rect 926 1858 930 1862
rect 974 1858 978 1862
rect 990 1858 994 1862
rect 1014 1858 1018 1862
rect 1046 1858 1050 1862
rect 1070 1858 1074 1862
rect 1118 1858 1122 1862
rect 1150 1858 1154 1862
rect 1174 1858 1178 1862
rect 1206 1858 1210 1862
rect 1222 1858 1226 1862
rect 1254 1858 1258 1862
rect 1286 1858 1290 1862
rect 1326 1858 1330 1862
rect 1350 1858 1354 1862
rect 1406 1858 1410 1862
rect 1462 1858 1466 1862
rect 1494 1858 1498 1862
rect 1526 1858 1530 1862
rect 1590 1858 1594 1862
rect 1622 1858 1626 1862
rect 1662 1858 1666 1862
rect 1670 1858 1674 1862
rect 1678 1858 1682 1862
rect 1702 1858 1706 1862
rect 1718 1858 1722 1862
rect 1750 1858 1754 1862
rect 1798 1858 1802 1862
rect 1910 1858 1914 1862
rect 1958 1858 1962 1862
rect 2038 1858 2042 1862
rect 2086 1858 2090 1862
rect 2102 1858 2106 1862
rect 2126 1858 2130 1862
rect 2134 1858 2138 1862
rect 2150 1858 2154 1862
rect 2174 1858 2178 1862
rect 2182 1858 2186 1862
rect 2206 1858 2210 1862
rect 2238 1858 2242 1862
rect 2294 1868 2298 1872
rect 2366 1868 2370 1872
rect 2430 1868 2434 1872
rect 2454 1868 2458 1872
rect 2502 1868 2506 1872
rect 2606 1868 2610 1872
rect 2694 1868 2698 1872
rect 2734 1868 2738 1872
rect 2798 1868 2802 1872
rect 2814 1868 2818 1872
rect 2950 1868 2954 1872
rect 2974 1868 2978 1872
rect 3078 1868 3082 1872
rect 3094 1868 3098 1872
rect 3110 1868 3114 1872
rect 3118 1868 3122 1872
rect 3142 1868 3146 1872
rect 2286 1858 2290 1862
rect 2310 1858 2314 1862
rect 2326 1858 2330 1862
rect 2334 1858 2338 1862
rect 2342 1858 2346 1862
rect 2406 1858 2410 1862
rect 2438 1858 2442 1862
rect 2470 1858 2474 1862
rect 2550 1858 2554 1862
rect 2678 1858 2682 1862
rect 2702 1858 2706 1862
rect 2726 1858 2730 1862
rect 2758 1858 2762 1862
rect 2790 1858 2794 1862
rect 2886 1858 2890 1862
rect 3046 1858 3050 1862
rect 3206 1868 3210 1872
rect 3214 1868 3218 1872
rect 3230 1868 3234 1872
rect 3246 1868 3250 1872
rect 3086 1858 3090 1862
rect 3102 1858 3106 1862
rect 3118 1858 3122 1862
rect 3158 1858 3162 1862
rect 3182 1858 3186 1862
rect 3198 1858 3202 1862
rect 3222 1858 3226 1862
rect 3270 1858 3274 1862
rect 3294 1858 3298 1862
rect 3310 1868 3314 1872
rect 3430 1868 3434 1872
rect 3526 1868 3530 1872
rect 3542 1868 3546 1872
rect 3558 1868 3562 1872
rect 3590 1868 3594 1872
rect 3638 1868 3642 1872
rect 3662 1868 3666 1872
rect 3678 1868 3682 1872
rect 3686 1868 3690 1872
rect 3718 1868 3722 1872
rect 3742 1868 3746 1872
rect 3758 1868 3762 1872
rect 3774 1868 3778 1872
rect 3790 1868 3794 1872
rect 3822 1868 3826 1872
rect 3894 1868 3898 1872
rect 4086 1868 4090 1872
rect 4246 1868 4250 1872
rect 4326 1868 4330 1872
rect 3374 1858 3378 1862
rect 3518 1858 3522 1862
rect 3550 1858 3554 1862
rect 3582 1858 3586 1862
rect 3598 1858 3602 1862
rect 3614 1858 3618 1862
rect 3646 1858 3650 1862
rect 3678 1858 3682 1862
rect 3686 1858 3690 1862
rect 3734 1858 3738 1862
rect 3766 1858 3770 1862
rect 3782 1858 3786 1862
rect 3830 1858 3834 1862
rect 3862 1858 3866 1862
rect 3910 1858 3914 1862
rect 3942 1858 3946 1862
rect 3966 1858 3970 1862
rect 3998 1858 4002 1862
rect 4022 1858 4026 1862
rect 4070 1858 4074 1862
rect 4118 1858 4122 1862
rect 4150 1858 4154 1862
rect 4190 1858 4194 1862
rect 4230 1858 4234 1862
rect 4294 1858 4298 1862
rect 4342 1858 4346 1862
rect 4350 1858 4354 1862
rect 4366 1858 4370 1862
rect 478 1848 482 1852
rect 486 1848 490 1852
rect 686 1848 690 1852
rect 702 1848 706 1852
rect 710 1848 714 1852
rect 798 1848 802 1852
rect 910 1848 914 1852
rect 958 1848 962 1852
rect 1030 1848 1034 1852
rect 1062 1848 1066 1852
rect 1134 1848 1138 1852
rect 1190 1848 1194 1852
rect 1222 1848 1226 1852
rect 1246 1848 1250 1852
rect 1302 1848 1306 1852
rect 1310 1848 1314 1852
rect 1366 1848 1370 1852
rect 1390 1848 1394 1852
rect 1446 1848 1450 1852
rect 1478 1848 1482 1852
rect 1550 1848 1554 1852
rect 1822 1850 1826 1854
rect 2054 1848 2058 1852
rect 2158 1848 2162 1852
rect 2214 1848 2218 1852
rect 2302 1848 2306 1852
rect 2310 1848 2314 1852
rect 2382 1848 2386 1852
rect 2406 1848 2410 1852
rect 2654 1848 2658 1852
rect 2710 1848 2714 1852
rect 2774 1848 2778 1852
rect 2806 1848 2810 1852
rect 3174 1848 3178 1852
rect 3182 1848 3186 1852
rect 3238 1848 3242 1852
rect 3278 1848 3282 1852
rect 3326 1848 3330 1852
rect 3462 1850 3466 1854
rect 3654 1848 3658 1852
rect 3838 1848 3842 1852
rect 3902 1848 3906 1852
rect 3934 1848 3938 1852
rect 4006 1848 4010 1852
rect 4014 1848 4018 1852
rect 4110 1848 4114 1852
rect 4142 1848 4146 1852
rect 4198 1848 4202 1852
rect 4334 1848 4338 1852
rect 6 1838 10 1842
rect 694 1838 698 1842
rect 782 1838 786 1842
rect 1126 1838 1130 1842
rect 1262 1838 1266 1842
rect 1414 1838 1418 1842
rect 2198 1838 2202 1842
rect 3334 1838 3338 1842
rect 3918 1838 3922 1842
rect 3950 1838 3954 1842
rect 3990 1838 3994 1842
rect 4030 1838 4034 1842
rect 4126 1838 4130 1842
rect 4142 1838 4146 1842
rect 4158 1838 4162 1842
rect 4166 1838 4170 1842
rect 4182 1838 4186 1842
rect 1102 1828 1106 1832
rect 1254 1828 1258 1832
rect 1822 1827 1826 1831
rect 3462 1827 3466 1831
rect 4262 1828 4266 1832
rect 238 1818 242 1822
rect 414 1818 418 1822
rect 486 1818 490 1822
rect 742 1818 746 1822
rect 1014 1818 1018 1822
rect 1350 1818 1354 1822
rect 1406 1818 1410 1822
rect 1734 1818 1738 1822
rect 1950 1818 1954 1822
rect 2190 1818 2194 1822
rect 2510 1818 2514 1822
rect 2654 1818 2658 1822
rect 3030 1818 3034 1822
rect 3726 1818 3730 1822
rect 3758 1818 3762 1822
rect 3862 1818 3866 1822
rect 3926 1818 3930 1822
rect 4038 1818 4042 1822
rect 4054 1818 4058 1822
rect 4070 1818 4074 1822
rect 4190 1818 4194 1822
rect 4214 1818 4218 1822
rect 4302 1818 4306 1822
rect 4318 1818 4322 1822
rect 394 1803 398 1807
rect 401 1803 405 1807
rect 1418 1803 1422 1807
rect 1425 1803 1429 1807
rect 2442 1803 2446 1807
rect 2449 1803 2453 1807
rect 3474 1803 3478 1807
rect 3481 1803 3485 1807
rect 206 1788 210 1792
rect 238 1788 242 1792
rect 462 1788 466 1792
rect 606 1788 610 1792
rect 646 1788 650 1792
rect 998 1788 1002 1792
rect 1110 1788 1114 1792
rect 1198 1788 1202 1792
rect 1222 1788 1226 1792
rect 1278 1788 1282 1792
rect 1318 1788 1322 1792
rect 1470 1788 1474 1792
rect 1566 1788 1570 1792
rect 1630 1788 1634 1792
rect 1654 1788 1658 1792
rect 1718 1788 1722 1792
rect 1934 1788 1938 1792
rect 2422 1788 2426 1792
rect 2846 1788 2850 1792
rect 2878 1788 2882 1792
rect 3118 1788 3122 1792
rect 3742 1788 3746 1792
rect 3758 1788 3762 1792
rect 3774 1788 3778 1792
rect 3990 1788 3994 1792
rect 4030 1788 4034 1792
rect 4094 1788 4098 1792
rect 4182 1788 4186 1792
rect 4246 1788 4250 1792
rect 4286 1788 4290 1792
rect 4310 1788 4314 1792
rect 366 1779 370 1783
rect 1606 1778 1610 1782
rect 1742 1778 1746 1782
rect 1982 1778 1986 1782
rect 3046 1779 3050 1783
rect 3262 1778 3266 1782
rect 3926 1779 3930 1783
rect 30 1768 34 1772
rect 958 1768 962 1772
rect 1102 1768 1106 1772
rect 1190 1768 1194 1772
rect 1230 1768 1234 1772
rect 1310 1768 1314 1772
rect 1438 1768 1442 1772
rect 2270 1768 2274 1772
rect 3358 1768 3362 1772
rect 3606 1768 3610 1772
rect 3998 1768 4002 1772
rect 4022 1768 4026 1772
rect 4062 1768 4066 1772
rect 4086 1768 4090 1772
rect 4126 1768 4130 1772
rect 4134 1768 4138 1772
rect 4150 1768 4154 1772
rect 4166 1768 4170 1772
rect 4190 1768 4194 1772
rect 4278 1768 4282 1772
rect 4318 1768 4322 1772
rect 206 1758 210 1762
rect 366 1756 370 1760
rect 430 1758 434 1762
rect 446 1758 450 1762
rect 606 1758 610 1762
rect 646 1758 650 1762
rect 798 1758 802 1762
rect 1078 1758 1082 1762
rect 1134 1758 1138 1762
rect 1206 1758 1210 1762
rect 1262 1758 1266 1762
rect 1294 1758 1298 1762
rect 1446 1758 1450 1762
rect 1510 1758 1514 1762
rect 1726 1758 1730 1762
rect 1774 1758 1778 1762
rect 1934 1758 1938 1762
rect 2014 1758 2018 1762
rect 2070 1758 2074 1762
rect 2086 1758 2090 1762
rect 2142 1758 2146 1762
rect 2158 1758 2162 1762
rect 2182 1758 2186 1762
rect 2214 1758 2218 1762
rect 2246 1758 2250 1762
rect 2422 1758 2426 1762
rect 2462 1758 2466 1762
rect 2478 1758 2482 1762
rect 22 1748 26 1752
rect 190 1748 194 1752
rect 206 1748 210 1752
rect 382 1748 386 1752
rect 430 1748 434 1752
rect 590 1748 594 1752
rect 606 1748 610 1752
rect 654 1748 658 1752
rect 830 1748 834 1752
rect 846 1748 850 1752
rect 886 1748 890 1752
rect 918 1748 922 1752
rect 934 1748 938 1752
rect 942 1748 946 1752
rect 1022 1748 1026 1752
rect 1046 1748 1050 1752
rect 1054 1748 1058 1752
rect 1094 1748 1098 1752
rect 1118 1748 1122 1752
rect 1150 1748 1154 1752
rect 1174 1748 1178 1752
rect 1198 1748 1202 1752
rect 1278 1748 1282 1752
rect 1302 1748 1306 1752
rect 1334 1748 1338 1752
rect 1350 1748 1354 1752
rect 1390 1748 1394 1752
rect 1398 1748 1402 1752
rect 1454 1748 1458 1752
rect 1478 1748 1482 1752
rect 1534 1748 1538 1752
rect 1550 1748 1554 1752
rect 1590 1748 1594 1752
rect 1614 1748 1618 1752
rect 1654 1748 1658 1752
rect 1670 1748 1674 1752
rect 1686 1748 1690 1752
rect 1774 1748 1778 1752
rect 1918 1748 1922 1752
rect 1998 1748 2002 1752
rect 2030 1748 2034 1752
rect 2046 1748 2050 1752
rect 2070 1748 2074 1752
rect 2086 1748 2090 1752
rect 2110 1748 2114 1752
rect 2190 1748 2194 1752
rect 2206 1748 2210 1752
rect 2230 1748 2234 1752
rect 2318 1748 2322 1752
rect 2414 1748 2418 1752
rect 2478 1748 2482 1752
rect 2526 1748 2530 1752
rect 2534 1748 2538 1752
rect 2590 1758 2594 1762
rect 2686 1758 2690 1762
rect 2798 1758 2802 1762
rect 2830 1758 2834 1762
rect 2862 1758 2866 1762
rect 3046 1756 3050 1760
rect 3110 1758 3114 1762
rect 2606 1748 2610 1752
rect 2646 1748 2650 1752
rect 2654 1748 2658 1752
rect 2702 1748 2706 1752
rect 2734 1748 2738 1752
rect 6 1738 10 1742
rect 158 1738 162 1742
rect 334 1738 338 1742
rect 422 1738 426 1742
rect 558 1738 562 1742
rect 694 1738 698 1742
rect 822 1738 826 1742
rect 838 1738 842 1742
rect 862 1738 866 1742
rect 910 1738 914 1742
rect 950 1738 954 1742
rect 1030 1738 1034 1742
rect 1054 1738 1058 1742
rect 2782 1748 2786 1752
rect 2814 1748 2818 1752
rect 2830 1748 2834 1752
rect 2878 1748 2882 1752
rect 3054 1748 3058 1752
rect 3094 1748 3098 1752
rect 3118 1748 3122 1752
rect 3150 1748 3154 1752
rect 3246 1758 3250 1762
rect 3302 1758 3306 1762
rect 3374 1758 3378 1762
rect 3622 1758 3626 1762
rect 3638 1758 3642 1762
rect 3646 1758 3650 1762
rect 3702 1758 3706 1762
rect 3182 1748 3186 1752
rect 3198 1748 3202 1752
rect 3238 1748 3242 1752
rect 3262 1748 3266 1752
rect 3270 1748 3274 1752
rect 3286 1748 3290 1752
rect 3294 1748 3298 1752
rect 3926 1756 3930 1760
rect 3982 1758 3986 1762
rect 4038 1758 4042 1762
rect 4046 1758 4050 1762
rect 4102 1758 4106 1762
rect 4110 1758 4114 1762
rect 4166 1758 4170 1762
rect 4174 1758 4178 1762
rect 4294 1758 4298 1762
rect 4302 1758 4306 1762
rect 4342 1758 4346 1762
rect 3334 1748 3338 1752
rect 3366 1748 3370 1752
rect 3390 1748 3394 1752
rect 3398 1748 3402 1752
rect 3430 1748 3434 1752
rect 3454 1748 3458 1752
rect 3502 1748 3506 1752
rect 3510 1748 3514 1752
rect 3534 1748 3538 1752
rect 3582 1748 3586 1752
rect 3614 1748 3618 1752
rect 3622 1748 3626 1752
rect 3662 1748 3666 1752
rect 3686 1748 3690 1752
rect 3734 1748 3738 1752
rect 3934 1748 3938 1752
rect 3990 1748 3994 1752
rect 4022 1748 4026 1752
rect 4054 1748 4058 1752
rect 4094 1748 4098 1752
rect 4118 1748 4122 1752
rect 4158 1748 4162 1752
rect 4182 1748 4186 1752
rect 4206 1748 4210 1752
rect 4262 1748 4266 1752
rect 4278 1748 4282 1752
rect 4310 1748 4314 1752
rect 4358 1748 4362 1752
rect 4390 1748 4394 1752
rect 1214 1738 1218 1742
rect 1254 1738 1258 1742
rect 1286 1738 1290 1742
rect 1326 1738 1330 1742
rect 1358 1738 1362 1742
rect 1382 1738 1386 1742
rect 1414 1738 1418 1742
rect 1526 1738 1530 1742
rect 1542 1738 1546 1742
rect 1558 1738 1562 1742
rect 1582 1738 1586 1742
rect 1646 1738 1650 1742
rect 1678 1738 1682 1742
rect 1702 1738 1706 1742
rect 1758 1738 1762 1742
rect 1886 1738 1890 1742
rect 1990 1738 1994 1742
rect 2022 1738 2026 1742
rect 2054 1738 2058 1742
rect 2062 1738 2066 1742
rect 2142 1738 2146 1742
rect 2166 1738 2170 1742
rect 2190 1738 2194 1742
rect 2222 1738 2226 1742
rect 2254 1738 2258 1742
rect 2374 1738 2378 1742
rect 2550 1738 2554 1742
rect 2566 1738 2570 1742
rect 2614 1738 2618 1742
rect 2662 1738 2666 1742
rect 2710 1738 2714 1742
rect 2742 1738 2746 1742
rect 2750 1738 2754 1742
rect 2774 1738 2778 1742
rect 2790 1738 2794 1742
rect 2806 1738 2810 1742
rect 2838 1738 2842 1742
rect 2886 1738 2890 1742
rect 3014 1738 3018 1742
rect 3086 1738 3090 1742
rect 3142 1738 3146 1742
rect 3166 1738 3170 1742
rect 3174 1738 3178 1742
rect 3190 1738 3194 1742
rect 3230 1738 3234 1742
rect 3278 1738 3282 1742
rect 3310 1738 3314 1742
rect 3342 1738 3346 1742
rect 3406 1738 3410 1742
rect 3422 1738 3426 1742
rect 3462 1738 3466 1742
rect 3550 1738 3554 1742
rect 3614 1738 3618 1742
rect 3654 1738 3658 1742
rect 3678 1738 3682 1742
rect 3726 1738 3730 1742
rect 3750 1738 3754 1742
rect 3766 1738 3770 1742
rect 3782 1738 3786 1742
rect 3894 1738 3898 1742
rect 4214 1738 4218 1742
rect 142 1728 146 1732
rect 318 1728 322 1732
rect 542 1728 546 1732
rect 710 1728 714 1732
rect 1366 1728 1370 1732
rect 1518 1728 1522 1732
rect 1566 1728 1570 1732
rect 1598 1728 1602 1732
rect 1702 1728 1706 1732
rect 1710 1728 1714 1732
rect 1734 1728 1738 1732
rect 1750 1728 1754 1732
rect 1870 1728 1874 1732
rect 1966 1728 1970 1732
rect 2014 1728 2018 1732
rect 2094 1728 2098 1732
rect 2134 1728 2138 1732
rect 2358 1728 2362 1732
rect 2502 1728 2506 1732
rect 2718 1728 2722 1732
rect 2766 1728 2770 1732
rect 2854 1728 2858 1732
rect 2998 1728 3002 1732
rect 3118 1728 3122 1732
rect 3134 1728 3138 1732
rect 3214 1728 3218 1732
rect 3350 1728 3354 1732
rect 3406 1728 3410 1732
rect 3438 1728 3442 1732
rect 3590 1728 3594 1732
rect 3878 1728 3882 1732
rect 4158 1728 4162 1732
rect 4230 1728 4234 1732
rect 462 1718 466 1722
rect 814 1718 818 1722
rect 870 1718 874 1722
rect 918 1718 922 1722
rect 1246 1718 1250 1722
rect 1334 1718 1338 1722
rect 1374 1718 1378 1722
rect 1494 1718 1498 1722
rect 1790 1718 1794 1722
rect 2030 1718 2034 1722
rect 2126 1718 2130 1722
rect 2174 1718 2178 1722
rect 2246 1718 2250 1722
rect 2278 1718 2282 1722
rect 2630 1718 2634 1722
rect 2670 1718 2674 1722
rect 2758 1718 2762 1722
rect 2918 1718 2922 1722
rect 3334 1718 3338 1722
rect 3374 1718 3378 1722
rect 3542 1718 3546 1722
rect 3566 1718 3570 1722
rect 3718 1718 3722 1722
rect 4054 1718 4058 1722
rect 4222 1718 4226 1722
rect 4246 1718 4250 1722
rect 4374 1718 4378 1722
rect 898 1703 902 1707
rect 905 1703 909 1707
rect 1930 1703 1934 1707
rect 1937 1703 1941 1707
rect 2954 1703 2958 1707
rect 2961 1703 2965 1707
rect 3978 1703 3982 1707
rect 3985 1703 3989 1707
rect 30 1688 34 1692
rect 270 1688 274 1692
rect 702 1688 706 1692
rect 830 1688 834 1692
rect 862 1688 866 1692
rect 974 1688 978 1692
rect 1038 1688 1042 1692
rect 1062 1688 1066 1692
rect 1070 1688 1074 1692
rect 1166 1688 1170 1692
rect 1230 1688 1234 1692
rect 1262 1688 1266 1692
rect 1294 1688 1298 1692
rect 1334 1688 1338 1692
rect 1494 1688 1498 1692
rect 1830 1688 1834 1692
rect 1846 1688 1850 1692
rect 1910 1688 1914 1692
rect 1958 1688 1962 1692
rect 1990 1688 1994 1692
rect 2102 1688 2106 1692
rect 2118 1688 2122 1692
rect 2582 1688 2586 1692
rect 2702 1688 2706 1692
rect 2862 1688 2866 1692
rect 2974 1688 2978 1692
rect 3166 1688 3170 1692
rect 3198 1688 3202 1692
rect 3438 1688 3442 1692
rect 3542 1688 3546 1692
rect 3630 1688 3634 1692
rect 3686 1688 3690 1692
rect 4022 1688 4026 1692
rect 4238 1688 4242 1692
rect 142 1678 146 1682
rect 502 1678 506 1682
rect 590 1678 594 1682
rect 1102 1678 1106 1682
rect 1182 1678 1186 1682
rect 1302 1678 1306 1682
rect 1310 1678 1314 1682
rect 1414 1678 1418 1682
rect 1438 1678 1442 1682
rect 1582 1678 1586 1682
rect 1590 1678 1594 1682
rect 1726 1678 1730 1682
rect 1742 1678 1746 1682
rect 1862 1678 1866 1682
rect 1878 1678 1882 1682
rect 2086 1678 2090 1682
rect 2262 1678 2266 1682
rect 2390 1678 2394 1682
rect 2486 1678 2490 1682
rect 2574 1678 2578 1682
rect 2694 1678 2698 1682
rect 2782 1678 2786 1682
rect 2830 1678 2834 1682
rect 3070 1678 3074 1682
rect 3294 1678 3298 1682
rect 6 1668 10 1672
rect 158 1668 162 1672
rect 246 1668 250 1672
rect 326 1668 330 1672
rect 334 1668 338 1672
rect 366 1668 370 1672
rect 382 1668 386 1672
rect 398 1668 402 1672
rect 478 1668 482 1672
rect 486 1668 490 1672
rect 606 1668 610 1672
rect 678 1668 682 1672
rect 774 1668 778 1672
rect 806 1668 810 1672
rect 838 1668 842 1672
rect 942 1668 946 1672
rect 950 1668 954 1672
rect 1014 1668 1018 1672
rect 1046 1668 1050 1672
rect 1094 1668 1098 1672
rect 1142 1668 1146 1672
rect 1206 1668 1210 1672
rect 1222 1668 1226 1672
rect 1254 1668 1258 1672
rect 1278 1668 1282 1672
rect 1350 1668 1354 1672
rect 1390 1668 1394 1672
rect 1422 1668 1426 1672
rect 1462 1668 1466 1672
rect 1542 1668 1546 1672
rect 1558 1668 1562 1672
rect 1574 1668 1578 1672
rect 1598 1668 1602 1672
rect 1630 1668 1634 1672
rect 1662 1668 1666 1672
rect 1670 1668 1674 1672
rect 1822 1668 1826 1672
rect 1838 1668 1842 1672
rect 1886 1668 1890 1672
rect 1918 1668 1922 1672
rect 1974 1668 1978 1672
rect 2030 1668 2034 1672
rect 2038 1668 2042 1672
rect 2054 1668 2058 1672
rect 2062 1668 2066 1672
rect 2110 1668 2114 1672
rect 2134 1668 2138 1672
rect 2142 1668 2146 1672
rect 2158 1668 2162 1672
rect 2278 1668 2282 1672
rect 2350 1668 2354 1672
rect 2366 1668 2370 1672
rect 2502 1668 2506 1672
rect 2590 1668 2594 1672
rect 2622 1668 2626 1672
rect 2654 1668 2658 1672
rect 2686 1668 2690 1672
rect 2742 1668 2746 1672
rect 2750 1668 2754 1672
rect 2814 1668 2818 1672
rect 2870 1668 2874 1672
rect 2942 1668 2946 1672
rect 2966 1668 2970 1672
rect 3086 1668 3090 1672
rect 3158 1668 3162 1672
rect 3206 1668 3210 1672
rect 3310 1668 3314 1672
rect 3414 1668 3418 1672
rect 3446 1668 3450 1672
rect 3598 1678 3602 1682
rect 3750 1678 3754 1682
rect 3830 1678 3834 1682
rect 4246 1678 4250 1682
rect 4318 1678 4322 1682
rect 3526 1668 3530 1672
rect 3534 1668 3538 1672
rect 3550 1668 3554 1672
rect 3558 1668 3562 1672
rect 3614 1668 3618 1672
rect 3630 1668 3634 1672
rect 3646 1668 3650 1672
rect 3654 1668 3658 1672
rect 3694 1668 3698 1672
rect 3702 1668 3706 1672
rect 3734 1668 3738 1672
rect 3846 1668 3850 1672
rect 4078 1668 4082 1672
rect 4222 1668 4226 1672
rect 4318 1668 4322 1672
rect 4334 1668 4338 1672
rect 4350 1668 4354 1672
rect 22 1658 26 1662
rect 206 1658 210 1662
rect 230 1658 234 1662
rect 358 1658 362 1662
rect 374 1658 378 1662
rect 606 1658 610 1662
rect 654 1658 658 1662
rect 686 1658 690 1662
rect 718 1658 722 1662
rect 750 1658 754 1662
rect 782 1658 786 1662
rect 790 1658 794 1662
rect 814 1658 818 1662
rect 846 1658 850 1662
rect 886 1658 890 1662
rect 910 1658 914 1662
rect 934 1658 938 1662
rect 950 1658 954 1662
rect 982 1658 986 1662
rect 1006 1658 1010 1662
rect 1022 1658 1026 1662
rect 1086 1658 1090 1662
rect 1118 1658 1122 1662
rect 1150 1658 1154 1662
rect 1206 1658 1210 1662
rect 1246 1658 1250 1662
rect 1278 1658 1282 1662
rect 1334 1658 1338 1662
rect 1358 1658 1362 1662
rect 1382 1658 1386 1662
rect 1398 1658 1402 1662
rect 1414 1658 1418 1662
rect 1438 1658 1442 1662
rect 1470 1658 1474 1662
rect 1478 1658 1482 1662
rect 1510 1658 1514 1662
rect 1534 1658 1538 1662
rect 1550 1658 1554 1662
rect 1566 1658 1570 1662
rect 1606 1658 1610 1662
rect 1622 1658 1626 1662
rect 1638 1658 1642 1662
rect 1654 1658 1658 1662
rect 1710 1658 1714 1662
rect 1734 1658 1738 1662
rect 1758 1658 1762 1662
rect 1790 1658 1794 1662
rect 1814 1658 1818 1662
rect 1862 1658 1866 1662
rect 1910 1658 1914 1662
rect 1942 1658 1946 1662
rect 2014 1658 2018 1662
rect 2030 1658 2034 1662
rect 2070 1658 2074 1662
rect 2150 1658 2154 1662
rect 2318 1658 2322 1662
rect 2405 1658 2409 1662
rect 2542 1658 2546 1662
rect 2598 1658 2602 1662
rect 2614 1658 2618 1662
rect 2638 1658 2642 1662
rect 2678 1658 2682 1662
rect 2710 1658 2714 1662
rect 2726 1658 2730 1662
rect 2734 1658 2738 1662
rect 2750 1658 2754 1662
rect 2766 1658 2770 1662
rect 2806 1658 2810 1662
rect 2846 1658 2850 1662
rect 3030 1658 3034 1662
rect 3126 1658 3130 1662
rect 3182 1658 3186 1662
rect 3254 1658 3258 1662
rect 3382 1658 3386 1662
rect 3414 1658 3418 1662
rect 3454 1658 3458 1662
rect 3494 1658 3498 1662
rect 3526 1658 3530 1662
rect 3566 1658 3570 1662
rect 3574 1658 3578 1662
rect 3622 1658 3626 1662
rect 3662 1658 3666 1662
rect 3710 1658 3714 1662
rect 3726 1658 3730 1662
rect 3886 1658 3890 1662
rect 3926 1658 3930 1662
rect 3958 1658 3962 1662
rect 4006 1658 4010 1662
rect 4038 1658 4042 1662
rect 4078 1658 4082 1662
rect 4102 1658 4106 1662
rect 4134 1658 4138 1662
rect 4166 1658 4170 1662
rect 4182 1658 4186 1662
rect 4198 1658 4202 1662
rect 4222 1658 4226 1662
rect 4262 1658 4266 1662
rect 4294 1658 4298 1662
rect 4342 1658 4346 1662
rect 4350 1658 4354 1662
rect 206 1648 210 1652
rect 390 1648 394 1652
rect 502 1648 506 1652
rect 638 1650 642 1654
rect 710 1648 714 1652
rect 742 1648 746 1652
rect 798 1648 802 1652
rect 830 1648 834 1652
rect 894 1648 898 1652
rect 918 1648 922 1652
rect 974 1648 978 1652
rect 1038 1648 1042 1652
rect 1070 1648 1074 1652
rect 1230 1648 1234 1652
rect 1262 1648 1266 1652
rect 1606 1648 1610 1652
rect 1638 1648 1642 1652
rect 1798 1648 1802 1652
rect 1814 1648 1818 1652
rect 1998 1648 2002 1652
rect 2094 1648 2098 1652
rect 2118 1648 2122 1652
rect 2174 1648 2178 1652
rect 2310 1650 2314 1654
rect 2550 1648 2554 1652
rect 2598 1648 2602 1652
rect 2630 1648 2634 1652
rect 2662 1648 2666 1652
rect 2718 1648 2722 1652
rect 2822 1648 2826 1652
rect 2830 1648 2834 1652
rect 3118 1650 3122 1654
rect 3198 1648 3202 1652
rect 3342 1650 3346 1654
rect 3438 1648 3442 1652
rect 3470 1648 3474 1652
rect 3518 1648 3522 1652
rect 3574 1648 3578 1652
rect 3630 1648 3634 1652
rect 3678 1648 3682 1652
rect 3726 1648 3730 1652
rect 3878 1650 3882 1654
rect 3918 1648 3922 1652
rect 3950 1648 3954 1652
rect 3998 1648 4002 1652
rect 4006 1648 4010 1652
rect 4030 1648 4034 1652
rect 4086 1648 4090 1652
rect 4094 1648 4098 1652
rect 4126 1648 4130 1652
rect 4158 1648 4162 1652
rect 4190 1648 4194 1652
rect 4254 1648 4258 1652
rect 4286 1648 4290 1652
rect 4358 1648 4362 1652
rect 4374 1648 4378 1652
rect 726 1638 730 1642
rect 758 1638 762 1642
rect 878 1638 882 1642
rect 1062 1638 1066 1642
rect 1774 1638 1778 1642
rect 2070 1638 2074 1642
rect 2174 1638 2178 1642
rect 3662 1638 3666 1642
rect 3934 1638 3938 1642
rect 3966 1638 3970 1642
rect 4014 1638 4018 1642
rect 4046 1638 4050 1642
rect 4070 1638 4074 1642
rect 4110 1638 4114 1642
rect 4142 1638 4146 1642
rect 4174 1638 4178 1642
rect 4198 1638 4202 1642
rect 4270 1638 4274 1642
rect 4294 1638 4298 1642
rect 1958 1628 1962 1632
rect 2310 1627 2314 1631
rect 3342 1627 3346 1631
rect 4214 1628 4218 1632
rect 206 1618 210 1622
rect 638 1618 642 1622
rect 750 1618 754 1622
rect 1134 1618 1138 1622
rect 1678 1618 1682 1622
rect 2054 1618 2058 1622
rect 2358 1618 2362 1622
rect 2550 1618 2554 1622
rect 2886 1618 2890 1622
rect 2990 1618 2994 1622
rect 3118 1618 3122 1622
rect 3398 1618 3402 1622
rect 3878 1618 3882 1622
rect 3942 1618 3946 1622
rect 4038 1618 4042 1622
rect 4102 1618 4106 1622
rect 4134 1618 4138 1622
rect 4262 1618 4266 1622
rect 4294 1618 4298 1622
rect 394 1603 398 1607
rect 401 1603 405 1607
rect 1418 1603 1422 1607
rect 1425 1603 1429 1607
rect 2442 1603 2446 1607
rect 2449 1603 2453 1607
rect 3474 1603 3478 1607
rect 3481 1603 3485 1607
rect 6 1588 10 1592
rect 102 1588 106 1592
rect 374 1588 378 1592
rect 422 1588 426 1592
rect 478 1588 482 1592
rect 694 1588 698 1592
rect 758 1588 762 1592
rect 902 1588 906 1592
rect 1174 1588 1178 1592
rect 1238 1588 1242 1592
rect 1350 1588 1354 1592
rect 1414 1588 1418 1592
rect 1566 1588 1570 1592
rect 1622 1588 1626 1592
rect 1814 1588 1818 1592
rect 2014 1588 2018 1592
rect 2166 1588 2170 1592
rect 2534 1588 2538 1592
rect 2934 1588 2938 1592
rect 3134 1588 3138 1592
rect 3382 1588 3386 1592
rect 3502 1588 3506 1592
rect 3838 1588 3842 1592
rect 4038 1588 4042 1592
rect 4198 1588 4202 1592
rect 4262 1588 4266 1592
rect 4278 1588 4282 1592
rect 4318 1588 4322 1592
rect 4342 1588 4346 1592
rect 30 1578 34 1582
rect 1110 1578 1114 1582
rect 126 1568 130 1572
rect 230 1568 234 1572
rect 646 1568 650 1572
rect 766 1568 770 1572
rect 1070 1568 1074 1572
rect 1102 1568 1106 1572
rect 2470 1579 2474 1583
rect 3006 1579 3010 1583
rect 3326 1578 3330 1582
rect 3438 1578 3442 1582
rect 3574 1578 3578 1582
rect 3646 1578 3650 1582
rect 1166 1568 1170 1572
rect 1198 1568 1202 1572
rect 1534 1568 1538 1572
rect 1598 1568 1602 1572
rect 1982 1568 1986 1572
rect 2070 1568 2074 1572
rect 2190 1568 2194 1572
rect 2262 1568 2266 1572
rect 3950 1568 3954 1572
rect 4030 1568 4034 1572
rect 4046 1568 4050 1572
rect 4062 1568 4066 1572
rect 4118 1568 4122 1572
rect 4150 1568 4154 1572
rect 4190 1568 4194 1572
rect 4222 1568 4226 1572
rect 4254 1568 4258 1572
rect 4286 1568 4290 1572
rect 4310 1568 4314 1572
rect 4350 1568 4354 1572
rect 62 1558 66 1562
rect 78 1558 82 1562
rect 142 1558 146 1562
rect 374 1558 378 1562
rect 478 1558 482 1562
rect 662 1558 666 1562
rect 710 1558 714 1562
rect 726 1558 730 1562
rect 750 1558 754 1562
rect 814 1558 818 1562
rect 846 1558 850 1562
rect 1054 1558 1058 1562
rect 1078 1558 1082 1562
rect 1086 1558 1090 1562
rect 1150 1558 1154 1562
rect 1182 1558 1186 1562
rect 1294 1558 1298 1562
rect 1470 1558 1474 1562
rect 1582 1558 1586 1562
rect 1614 1558 1618 1562
rect 1638 1558 1642 1562
rect 1694 1558 1698 1562
rect 1726 1558 1730 1562
rect 1774 1558 1778 1562
rect 1830 1558 1834 1562
rect 1838 1558 1842 1562
rect 1926 1558 1930 1562
rect 1966 1558 1970 1562
rect 1998 1558 2002 1562
rect 2150 1558 2154 1562
rect 2182 1558 2186 1562
rect 2230 1558 2234 1562
rect 22 1548 26 1552
rect 54 1548 58 1552
rect 62 1548 66 1552
rect 78 1548 82 1552
rect 126 1548 130 1552
rect 270 1548 274 1552
rect 382 1548 386 1552
rect 454 1548 458 1552
rect 478 1548 482 1552
rect 582 1548 586 1552
rect 638 1548 642 1552
rect 670 1548 674 1552
rect 694 1548 698 1552
rect 742 1548 746 1552
rect 758 1548 762 1552
rect 782 1548 786 1552
rect 830 1548 834 1552
rect 862 1548 866 1552
rect 886 1548 890 1552
rect 902 1548 906 1552
rect 942 1548 946 1552
rect 958 1548 962 1552
rect 1030 1548 1034 1552
rect 1062 1548 1066 1552
rect 1094 1548 1098 1552
rect 1126 1548 1130 1552
rect 1158 1548 1162 1552
rect 1190 1548 1194 1552
rect 54 1538 58 1542
rect 150 1538 154 1542
rect 214 1538 218 1542
rect 326 1538 330 1542
rect 398 1538 402 1542
rect 430 1538 434 1542
rect 526 1538 530 1542
rect 623 1538 627 1542
rect 630 1538 634 1542
rect 1270 1548 1274 1552
rect 1294 1548 1298 1552
rect 1310 1548 1314 1552
rect 1326 1548 1330 1552
rect 1366 1548 1370 1552
rect 1454 1548 1458 1552
rect 1510 1548 1514 1552
rect 1518 1548 1522 1552
rect 1542 1548 1546 1552
rect 1550 1548 1554 1552
rect 1566 1548 1570 1552
rect 1590 1548 1594 1552
rect 1654 1548 1658 1552
rect 1678 1548 1682 1552
rect 1710 1548 1714 1552
rect 1734 1548 1738 1552
rect 1750 1548 1754 1552
rect 1790 1548 1794 1552
rect 1814 1548 1818 1552
rect 1862 1548 1866 1552
rect 1894 1548 1898 1552
rect 1910 1548 1914 1552
rect 1950 1548 1954 1552
rect 2022 1548 2026 1552
rect 2054 1548 2058 1552
rect 2062 1548 2066 1552
rect 2070 1548 2074 1552
rect 2126 1548 2130 1552
rect 2134 1548 2138 1552
rect 2214 1548 2218 1552
rect 2302 1558 2306 1562
rect 2254 1548 2258 1552
rect 2286 1548 2290 1552
rect 2470 1556 2474 1560
rect 2598 1558 2602 1562
rect 2614 1558 2618 1562
rect 2718 1558 2722 1562
rect 2934 1558 2938 1562
rect 2942 1558 2946 1562
rect 2486 1548 2490 1552
rect 2550 1548 2554 1552
rect 2566 1548 2570 1552
rect 2590 1548 2594 1552
rect 2598 1548 2602 1552
rect 2622 1548 2626 1552
rect 2638 1548 2642 1552
rect 686 1538 690 1542
rect 782 1538 786 1542
rect 814 1538 818 1542
rect 838 1538 842 1542
rect 870 1538 874 1542
rect 878 1538 882 1542
rect 918 1538 922 1542
rect 950 1538 954 1542
rect 966 1538 970 1542
rect 974 1538 978 1542
rect 1006 1538 1010 1542
rect 1038 1538 1042 1542
rect 1118 1538 1122 1542
rect 1214 1538 1218 1542
rect 1254 1538 1258 1542
rect 1262 1538 1266 1542
rect 1286 1538 1290 1542
rect 1318 1538 1322 1542
rect 1334 1538 1338 1542
rect 1358 1538 1362 1542
rect 1390 1538 1394 1542
rect 1446 1538 1450 1542
rect 1478 1538 1482 1542
rect 1558 1538 1562 1542
rect 1590 1538 1594 1542
rect 1662 1538 1666 1542
rect 1686 1538 1690 1542
rect 1702 1538 1706 1542
rect 1734 1538 1738 1542
rect 1742 1538 1746 1542
rect 1798 1538 1802 1542
rect 1806 1538 1810 1542
rect 1862 1538 1866 1542
rect 1870 1538 1874 1542
rect 1902 1538 1906 1542
rect 1950 1538 1954 1542
rect 1974 1538 1978 1542
rect 2094 1538 2098 1542
rect 2102 1540 2106 1544
rect 2678 1548 2682 1552
rect 2710 1548 2714 1552
rect 2734 1548 2738 1552
rect 2750 1548 2754 1552
rect 2830 1548 2834 1552
rect 3006 1556 3010 1560
rect 3302 1558 3306 1562
rect 3310 1558 3314 1562
rect 3342 1558 3346 1562
rect 3470 1558 3474 1562
rect 3614 1558 3618 1562
rect 3630 1558 3634 1562
rect 3686 1558 3690 1562
rect 3694 1558 3698 1562
rect 3862 1558 3866 1562
rect 3934 1558 3938 1562
rect 4014 1558 4018 1562
rect 4046 1558 4050 1562
rect 4134 1558 4138 1562
rect 4166 1558 4170 1562
rect 4174 1558 4178 1562
rect 4206 1558 4210 1562
rect 4238 1558 4242 1562
rect 4270 1558 4274 1562
rect 4326 1558 4330 1562
rect 4334 1558 4338 1562
rect 2990 1548 2994 1552
rect 3174 1548 3178 1552
rect 3182 1548 3186 1552
rect 3246 1548 3250 1552
rect 3270 1548 3274 1552
rect 3286 1548 3290 1552
rect 3334 1548 3338 1552
rect 3366 1548 3370 1552
rect 3382 1548 3386 1552
rect 3398 1548 3402 1552
rect 3414 1548 3418 1552
rect 3454 1548 3458 1552
rect 3494 1548 3498 1552
rect 3510 1548 3514 1552
rect 3542 1548 3546 1552
rect 3550 1548 3554 1552
rect 3582 1548 3586 1552
rect 3606 1548 3610 1552
rect 3630 1548 3634 1552
rect 3670 1548 3674 1552
rect 3718 1548 3722 1552
rect 3726 1548 3730 1552
rect 3766 1548 3770 1552
rect 3782 1548 3786 1552
rect 3814 1548 3818 1552
rect 3822 1548 3826 1552
rect 3846 1548 3850 1552
rect 3910 1548 3914 1552
rect 3942 1548 3946 1552
rect 4022 1548 4026 1552
rect 4054 1548 4058 1552
rect 4150 1548 4154 1552
rect 4182 1548 4186 1552
rect 4214 1548 4218 1552
rect 4246 1548 4250 1552
rect 4278 1548 4282 1552
rect 4318 1548 4322 1552
rect 4342 1548 4346 1552
rect 2126 1538 2130 1542
rect 2158 1538 2162 1542
rect 2254 1538 2258 1542
rect 2334 1538 2338 1542
rect 2438 1538 2442 1542
rect 2510 1538 2514 1542
rect 2558 1538 2562 1542
rect 2574 1538 2578 1542
rect 2590 1538 2594 1542
rect 2630 1538 2634 1542
rect 2654 1538 2658 1542
rect 2686 1538 2690 1542
rect 2742 1538 2746 1542
rect 2782 1538 2786 1542
rect 2886 1538 2890 1542
rect 3038 1538 3042 1542
rect 3150 1538 3154 1542
rect 3166 1538 3170 1542
rect 3214 1538 3218 1542
rect 3278 1538 3282 1542
rect 3334 1538 3338 1542
rect 3350 1538 3354 1542
rect 3366 1538 3370 1542
rect 3374 1538 3378 1542
rect 3406 1538 3410 1542
rect 3422 1538 3426 1542
rect 3438 1538 3442 1542
rect 3526 1538 3530 1542
rect 3558 1538 3562 1542
rect 3574 1538 3578 1542
rect 3654 1538 3658 1542
rect 3662 1538 3666 1542
rect 3702 1538 3706 1542
rect 3718 1538 3722 1542
rect 3726 1538 3730 1542
rect 3774 1538 3778 1542
rect 3790 1538 3794 1542
rect 3854 1538 3858 1542
rect 3902 1538 3906 1542
rect 3910 1538 3914 1542
rect 3926 1538 3930 1542
rect 3990 1538 3994 1542
rect 4006 1538 4010 1542
rect 4086 1538 4090 1542
rect 4110 1538 4114 1542
rect 4158 1538 4162 1542
rect 4230 1538 4234 1542
rect 310 1528 314 1532
rect 542 1528 546 1532
rect 1278 1528 1282 1532
rect 1350 1528 1354 1532
rect 1366 1528 1370 1532
rect 1414 1528 1418 1532
rect 1438 1528 1442 1532
rect 1630 1528 1634 1532
rect 2006 1528 2010 1532
rect 2086 1528 2090 1532
rect 2190 1528 2194 1532
rect 2262 1528 2266 1532
rect 2422 1528 2426 1532
rect 2646 1528 2650 1532
rect 2654 1528 2658 1532
rect 2686 1528 2690 1532
rect 2790 1528 2794 1532
rect 2870 1528 2874 1532
rect 3054 1528 3058 1532
rect 3158 1528 3162 1532
rect 3254 1528 3258 1532
rect 3302 1528 3306 1532
rect 3438 1528 3442 1532
rect 3510 1528 3514 1532
rect 3590 1528 3594 1532
rect 3686 1528 3690 1532
rect 3750 1528 3754 1532
rect 3798 1528 3802 1532
rect 3886 1528 3890 1532
rect 4006 1528 4010 1532
rect 4102 1528 4106 1532
rect 806 1518 810 1522
rect 846 1518 850 1522
rect 1014 1518 1018 1522
rect 1094 1518 1098 1522
rect 1142 1518 1146 1522
rect 1198 1518 1202 1522
rect 1222 1518 1226 1522
rect 1470 1518 1474 1522
rect 1638 1518 1642 1522
rect 1766 1518 1770 1522
rect 1774 1518 1778 1522
rect 1838 1518 1842 1522
rect 2038 1518 2042 1522
rect 2318 1518 2322 1522
rect 2342 1518 2346 1522
rect 2694 1518 2698 1522
rect 3222 1518 3226 1522
rect 3478 1518 3482 1522
rect 3502 1518 3506 1522
rect 3598 1518 3602 1522
rect 3806 1518 3810 1522
rect 3838 1518 3842 1522
rect 898 1503 902 1507
rect 905 1503 909 1507
rect 1930 1503 1934 1507
rect 1937 1503 1941 1507
rect 2954 1503 2958 1507
rect 2961 1503 2965 1507
rect 3978 1503 3982 1507
rect 3985 1503 3989 1507
rect 6 1488 10 1492
rect 270 1488 274 1492
rect 630 1488 634 1492
rect 702 1488 706 1492
rect 822 1488 826 1492
rect 854 1488 858 1492
rect 982 1488 986 1492
rect 1054 1488 1058 1492
rect 1262 1488 1266 1492
rect 1342 1488 1346 1492
rect 1366 1488 1370 1492
rect 1430 1488 1434 1492
rect 1462 1488 1466 1492
rect 1478 1488 1482 1492
rect 1502 1488 1506 1492
rect 1646 1488 1650 1492
rect 1902 1488 1906 1492
rect 2134 1488 2138 1492
rect 2374 1488 2378 1492
rect 2414 1488 2418 1492
rect 3102 1488 3106 1492
rect 3302 1488 3306 1492
rect 3422 1488 3426 1492
rect 3654 1488 3658 1492
rect 3678 1488 3682 1492
rect 3814 1488 3818 1492
rect 3846 1488 3850 1492
rect 4294 1488 4298 1492
rect 86 1478 90 1482
rect 166 1478 170 1482
rect 366 1478 370 1482
rect 486 1478 490 1482
rect 798 1478 802 1482
rect 878 1478 882 1482
rect 1166 1478 1170 1482
rect 1254 1478 1258 1482
rect 1398 1478 1402 1482
rect 1422 1478 1426 1482
rect 1486 1478 1490 1482
rect 1534 1478 1538 1482
rect 1622 1478 1626 1482
rect 1686 1478 1690 1482
rect 1718 1478 1722 1482
rect 1758 1478 1762 1482
rect 1766 1478 1770 1482
rect 1830 1478 1834 1482
rect 1846 1478 1850 1482
rect 1870 1478 1874 1482
rect 1934 1478 1938 1482
rect 2214 1478 2218 1482
rect 2566 1478 2570 1482
rect 2774 1478 2778 1482
rect 2782 1478 2786 1482
rect 2806 1478 2810 1482
rect 2830 1478 2834 1482
rect 2854 1478 2858 1482
rect 2982 1478 2986 1482
rect 3206 1478 3210 1482
rect 3310 1478 3314 1482
rect 3390 1478 3394 1482
rect 3454 1478 3458 1482
rect 3534 1478 3538 1482
rect 3590 1478 3594 1482
rect 3702 1478 3706 1482
rect 3742 1478 3746 1482
rect 3766 1478 3770 1482
rect 3774 1478 3778 1482
rect 3942 1478 3946 1482
rect 4166 1478 4170 1482
rect 4262 1478 4266 1482
rect 4310 1478 4314 1482
rect 54 1468 58 1472
rect 62 1468 66 1472
rect 182 1468 186 1472
rect 350 1468 354 1472
rect 470 1468 474 1472
rect 526 1468 530 1472
rect 654 1468 658 1472
rect 670 1468 674 1472
rect 718 1468 722 1472
rect 750 1468 754 1472
rect 838 1468 842 1472
rect 862 1468 866 1472
rect 910 1468 914 1472
rect 926 1468 930 1472
rect 934 1468 938 1472
rect 1014 1468 1018 1472
rect 1070 1468 1074 1472
rect 1182 1468 1186 1472
rect 1270 1468 1274 1472
rect 1318 1468 1322 1472
rect 1350 1468 1354 1472
rect 1358 1468 1362 1472
rect 1390 1468 1394 1472
rect 1446 1468 1450 1472
rect 1470 1468 1474 1472
rect 1494 1468 1498 1472
rect 1582 1468 1586 1472
rect 1614 1468 1618 1472
rect 1670 1468 1674 1472
rect 1678 1468 1682 1472
rect 1710 1468 1714 1472
rect 1806 1468 1810 1472
rect 1822 1468 1826 1472
rect 1878 1468 1882 1472
rect 1998 1468 2002 1472
rect 2030 1468 2034 1472
rect 2070 1468 2074 1472
rect 2230 1468 2234 1472
rect 2302 1468 2306 1472
rect 2334 1468 2338 1472
rect 2398 1468 2402 1472
rect 2422 1468 2426 1472
rect 2462 1468 2466 1472
rect 2485 1468 2489 1472
rect 2582 1468 2586 1472
rect 2654 1468 2658 1472
rect 2670 1468 2674 1472
rect 2686 1468 2690 1472
rect 2694 1468 2698 1472
rect 2718 1468 2722 1472
rect 2734 1468 2738 1472
rect 2758 1468 2762 1472
rect 2998 1468 3002 1472
rect 3110 1468 3114 1472
rect 3222 1468 3226 1472
rect 3318 1468 3322 1472
rect 3334 1468 3338 1472
rect 3350 1468 3354 1472
rect 3382 1468 3386 1472
rect 3406 1468 3410 1472
rect 3446 1468 3450 1472
rect 3558 1468 3562 1472
rect 3574 1468 3578 1472
rect 3606 1468 3610 1472
rect 3630 1468 3634 1472
rect 3790 1468 3794 1472
rect 3830 1468 3834 1472
rect 3958 1468 3962 1472
rect 4062 1468 4066 1472
rect 4166 1468 4170 1472
rect 4198 1468 4202 1472
rect 4246 1468 4250 1472
rect 54 1458 58 1462
rect 62 1458 66 1462
rect 78 1458 82 1462
rect 182 1458 186 1462
rect 254 1458 258 1462
rect 302 1458 306 1462
rect 478 1458 482 1462
rect 494 1458 498 1462
rect 510 1458 514 1462
rect 518 1458 522 1462
rect 566 1458 570 1462
rect 598 1458 602 1462
rect 646 1458 650 1462
rect 654 1458 658 1462
rect 686 1458 690 1462
rect 726 1458 730 1462
rect 742 1458 746 1462
rect 782 1458 786 1462
rect 814 1458 818 1462
rect 870 1458 874 1462
rect 878 1458 882 1462
rect 982 1458 986 1462
rect 1038 1458 1042 1462
rect 1126 1458 1130 1462
rect 1278 1458 1282 1462
rect 1286 1458 1290 1462
rect 1326 1458 1330 1462
rect 1342 1458 1346 1462
rect 1366 1458 1370 1462
rect 1382 1458 1386 1462
rect 1518 1458 1522 1462
rect 1566 1458 1570 1462
rect 1590 1458 1594 1462
rect 1598 1458 1602 1462
rect 1638 1458 1642 1462
rect 1662 1458 1666 1462
rect 1686 1458 1690 1462
rect 1742 1458 1746 1462
rect 1782 1458 1786 1462
rect 1798 1458 1802 1462
rect 1814 1458 1818 1462
rect 1830 1458 1834 1462
rect 1854 1458 1858 1462
rect 1902 1458 1906 1462
rect 1918 1458 1922 1462
rect 1958 1458 1962 1462
rect 1966 1458 1970 1462
rect 1990 1458 1994 1462
rect 2022 1458 2026 1462
rect 2038 1458 2042 1462
rect 2118 1458 2122 1462
rect 2270 1458 2274 1462
rect 2310 1458 2314 1462
rect 2326 1458 2330 1462
rect 2358 1458 2362 1462
rect 2398 1458 2402 1462
rect 2478 1458 2482 1462
rect 2526 1458 2530 1462
rect 2630 1458 2634 1462
rect 2654 1458 2658 1462
rect 2694 1458 2698 1462
rect 2726 1458 2730 1462
rect 2742 1458 2746 1462
rect 2766 1458 2770 1462
rect 2790 1458 2794 1462
rect 2798 1458 2802 1462
rect 2822 1458 2826 1462
rect 2846 1458 2850 1462
rect 2870 1458 2874 1462
rect 2901 1458 2905 1462
rect 3046 1458 3050 1462
rect 3086 1458 3090 1462
rect 3166 1458 3170 1462
rect 3270 1458 3274 1462
rect 3294 1458 3298 1462
rect 3326 1458 3330 1462
rect 3342 1458 3346 1462
rect 3358 1458 3362 1462
rect 3374 1458 3378 1462
rect 3414 1458 3418 1462
rect 3438 1458 3442 1462
rect 3470 1458 3474 1462
rect 3510 1458 3514 1462
rect 3550 1458 3554 1462
rect 3566 1458 3570 1462
rect 3622 1458 3626 1462
rect 3670 1458 3674 1462
rect 3694 1458 3698 1462
rect 3718 1458 3722 1462
rect 3726 1458 3730 1462
rect 3750 1458 3754 1462
rect 3790 1458 3794 1462
rect 3798 1458 3802 1462
rect 3902 1458 3906 1462
rect 4062 1458 4066 1462
rect 4086 1458 4090 1462
rect 4102 1458 4106 1462
rect 4118 1458 4122 1462
rect 4142 1458 4146 1462
rect 4182 1458 4186 1462
rect 4214 1458 4218 1462
rect 4238 1458 4242 1462
rect 4278 1458 4282 1462
rect 4326 1458 4330 1462
rect 4358 1458 4362 1462
rect 4390 1458 4394 1462
rect 30 1448 34 1452
rect 230 1448 234 1452
rect 302 1448 306 1452
rect 494 1448 498 1452
rect 550 1448 554 1452
rect 558 1448 562 1452
rect 590 1448 594 1452
rect 678 1448 682 1452
rect 846 1448 850 1452
rect 990 1448 994 1452
rect 1046 1448 1050 1452
rect 1054 1448 1058 1452
rect 1214 1450 1218 1454
rect 1406 1448 1410 1452
rect 1454 1448 1458 1452
rect 1646 1448 1650 1452
rect 2006 1448 2010 1452
rect 2054 1448 2058 1452
rect 2086 1448 2090 1452
rect 2110 1448 2114 1452
rect 2262 1450 2266 1454
rect 2326 1448 2330 1452
rect 2414 1448 2418 1452
rect 2438 1448 2442 1452
rect 2630 1448 2634 1452
rect 2710 1448 2714 1452
rect 2742 1448 2746 1452
rect 3046 1448 3050 1452
rect 3070 1448 3074 1452
rect 3086 1448 3090 1452
rect 3254 1450 3258 1454
rect 3358 1448 3362 1452
rect 3390 1448 3394 1452
rect 3422 1448 3426 1452
rect 3494 1448 3498 1452
rect 3582 1448 3586 1452
rect 3638 1448 3642 1452
rect 3678 1448 3682 1452
rect 3846 1448 3850 1452
rect 3990 1450 3994 1454
rect 4070 1448 4074 1452
rect 4078 1448 4082 1452
rect 4110 1448 4114 1452
rect 4174 1448 4178 1452
rect 4206 1448 4210 1452
rect 4294 1448 4298 1452
rect 574 1438 578 1442
rect 598 1438 602 1442
rect 606 1438 610 1442
rect 822 1438 826 1442
rect 886 1438 890 1442
rect 974 1438 978 1442
rect 1006 1438 1010 1442
rect 1030 1438 1034 1442
rect 1510 1438 1514 1442
rect 2022 1438 2026 1442
rect 4054 1438 4058 1442
rect 4094 1438 4098 1442
rect 4126 1438 4130 1442
rect 4190 1438 4194 1442
rect 4222 1438 4226 1442
rect 534 1428 538 1432
rect 566 1428 570 1432
rect 1214 1427 1218 1431
rect 2134 1428 2138 1432
rect 2262 1427 2266 1431
rect 4214 1428 4218 1432
rect 4342 1428 4346 1432
rect 230 1418 234 1422
rect 302 1418 306 1422
rect 726 1418 730 1422
rect 766 1418 770 1422
rect 830 1418 834 1422
rect 894 1418 898 1422
rect 982 1418 986 1422
rect 1038 1418 1042 1422
rect 1086 1418 1090 1422
rect 1302 1418 1306 1422
rect 1750 1418 1754 1422
rect 2430 1418 2434 1422
rect 2630 1418 2634 1422
rect 2814 1418 2818 1422
rect 2838 1418 2842 1422
rect 2878 1418 2882 1422
rect 3046 1418 3050 1422
rect 3254 1418 3258 1422
rect 3606 1418 3610 1422
rect 3734 1418 3738 1422
rect 3750 1418 3754 1422
rect 3814 1418 3818 1422
rect 3862 1418 3866 1422
rect 3990 1418 3994 1422
rect 4374 1418 4378 1422
rect 394 1403 398 1407
rect 401 1403 405 1407
rect 1418 1403 1422 1407
rect 1425 1403 1429 1407
rect 2442 1403 2446 1407
rect 2449 1403 2453 1407
rect 3474 1403 3478 1407
rect 3481 1403 3485 1407
rect 86 1388 90 1392
rect 294 1388 298 1392
rect 486 1388 490 1392
rect 526 1388 530 1392
rect 766 1388 770 1392
rect 862 1388 866 1392
rect 1206 1388 1210 1392
rect 1254 1388 1258 1392
rect 1326 1388 1330 1392
rect 1502 1388 1506 1392
rect 1558 1388 1562 1392
rect 1702 1388 1706 1392
rect 1902 1388 1906 1392
rect 2030 1388 2034 1392
rect 2070 1388 2074 1392
rect 2102 1388 2106 1392
rect 2262 1388 2266 1392
rect 3214 1388 3218 1392
rect 3270 1388 3274 1392
rect 3406 1388 3410 1392
rect 3590 1388 3594 1392
rect 3742 1388 3746 1392
rect 3910 1388 3914 1392
rect 3942 1388 3946 1392
rect 4054 1388 4058 1392
rect 4086 1388 4090 1392
rect 4102 1388 4106 1392
rect 4182 1388 4186 1392
rect 4238 1388 4242 1392
rect 4302 1388 4306 1392
rect 4326 1388 4330 1392
rect 150 1378 154 1382
rect 342 1378 346 1382
rect 1982 1378 1986 1382
rect 2118 1378 2122 1382
rect 2358 1378 2362 1382
rect 2494 1378 2498 1382
rect 6 1368 10 1372
rect 30 1368 34 1372
rect 62 1368 66 1372
rect 686 1368 690 1372
rect 798 1368 802 1372
rect 806 1368 810 1372
rect 862 1368 866 1372
rect 3694 1368 3698 1372
rect 3830 1368 3834 1372
rect 3902 1368 3906 1372
rect 3934 1368 3938 1372
rect 3966 1368 3970 1372
rect 4046 1368 4050 1372
rect 4078 1368 4082 1372
rect 4126 1368 4130 1372
rect 4142 1368 4146 1372
rect 4174 1368 4178 1372
rect 4230 1368 4234 1372
rect 4294 1368 4298 1372
rect 78 1358 82 1362
rect 118 1358 122 1362
rect 134 1358 138 1362
rect 294 1358 298 1362
rect 302 1358 306 1362
rect 486 1358 490 1362
rect 494 1358 498 1362
rect 526 1358 530 1362
rect 750 1358 754 1362
rect 782 1358 786 1362
rect 790 1358 794 1362
rect 822 1358 826 1362
rect 854 1358 858 1362
rect 894 1358 898 1362
rect 910 1358 914 1362
rect 942 1358 946 1362
rect 958 1358 962 1362
rect 1086 1358 1090 1362
rect 1222 1358 1226 1362
rect 1318 1358 1322 1362
rect 1414 1358 1418 1362
rect 1430 1358 1434 1362
rect 1478 1358 1482 1362
rect 1662 1358 1666 1362
rect 22 1348 26 1352
rect 46 1348 50 1352
rect 54 1348 58 1352
rect 102 1348 106 1352
rect 118 1348 122 1352
rect 190 1348 194 1352
rect 382 1348 386 1352
rect 526 1348 530 1352
rect 710 1348 714 1352
rect 734 1348 738 1352
rect 766 1348 770 1352
rect 798 1348 802 1352
rect 822 1348 826 1352
rect 838 1348 842 1352
rect 862 1348 866 1352
rect 894 1348 898 1352
rect 926 1348 930 1352
rect 1006 1348 1010 1352
rect 1046 1348 1050 1352
rect 1062 1348 1066 1352
rect 1102 1348 1106 1352
rect 1150 1348 1154 1352
rect 1158 1348 1162 1352
rect 1182 1348 1186 1352
rect 1238 1348 1242 1352
rect 1254 1348 1258 1352
rect 1294 1348 1298 1352
rect 1342 1348 1346 1352
rect 1350 1348 1354 1352
rect 1374 1348 1378 1352
rect 1462 1348 1466 1352
rect 1486 1348 1490 1352
rect 1590 1348 1594 1352
rect 1606 1348 1610 1352
rect 1654 1348 1658 1352
rect 1670 1348 1674 1352
rect 1686 1348 1690 1352
rect 1718 1358 1722 1362
rect 1838 1358 1842 1362
rect 1846 1358 1850 1362
rect 1862 1358 1866 1362
rect 1878 1358 1882 1362
rect 1926 1358 1930 1362
rect 2262 1358 2266 1362
rect 2294 1358 2298 1362
rect 2310 1358 2314 1362
rect 2342 1358 2346 1362
rect 2438 1358 2442 1362
rect 2590 1358 2594 1362
rect 2678 1358 2682 1362
rect 2734 1358 2738 1362
rect 2790 1358 2794 1362
rect 2814 1358 2818 1362
rect 2846 1358 2850 1362
rect 2966 1358 2970 1362
rect 2998 1358 3002 1362
rect 3214 1358 3218 1362
rect 3238 1358 3242 1362
rect 3318 1358 3322 1362
rect 3334 1358 3338 1362
rect 3366 1358 3370 1362
rect 3590 1358 3594 1362
rect 3614 1358 3618 1362
rect 3726 1358 3730 1362
rect 3790 1358 3794 1362
rect 3798 1358 3802 1362
rect 3886 1358 3890 1362
rect 3918 1358 3922 1362
rect 3950 1358 3954 1362
rect 4030 1358 4034 1362
rect 4062 1358 4066 1362
rect 4118 1358 4122 1362
rect 4158 1358 4162 1362
rect 4214 1358 4218 1362
rect 4246 1358 4250 1362
rect 4278 1358 4282 1362
rect 4310 1358 4314 1362
rect 4342 1358 4346 1362
rect 1734 1348 1738 1352
rect 1750 1348 1754 1352
rect 1774 1348 1778 1352
rect 1790 1348 1794 1352
rect 1822 1348 1826 1352
rect 1878 1348 1882 1352
rect 1902 1348 1906 1352
rect 1966 1348 1970 1352
rect 1990 1348 1994 1352
rect 2006 1348 2010 1352
rect 2022 1348 2026 1352
rect 2046 1348 2050 1352
rect 2054 1348 2058 1352
rect 2062 1348 2066 1352
rect 2102 1348 2106 1352
rect 2158 1348 2162 1352
rect 2270 1348 2274 1352
rect 2294 1348 2298 1352
rect 2326 1348 2330 1352
rect 2334 1348 2338 1352
rect 2382 1348 2386 1352
rect 2398 1348 2402 1352
rect 2430 1348 2434 1352
rect 2470 1348 2474 1352
rect 2502 1348 2506 1352
rect 2550 1348 2554 1352
rect 2566 1348 2570 1352
rect 2574 1348 2578 1352
rect 2598 1348 2602 1352
rect 2622 1348 2626 1352
rect 2630 1348 2634 1352
rect 2662 1348 2666 1352
rect 2678 1348 2682 1352
rect 2726 1348 2730 1352
rect 2782 1348 2786 1352
rect 2814 1348 2818 1352
rect 2830 1348 2834 1352
rect 2862 1348 2866 1352
rect 2878 1348 2882 1352
rect 2918 1348 2922 1352
rect 2966 1348 2970 1352
rect 3014 1348 3018 1352
rect 3054 1348 3058 1352
rect 3166 1348 3170 1352
rect 3262 1348 3266 1352
rect 3310 1348 3314 1352
rect 3334 1348 3338 1352
rect 3382 1348 3386 1352
rect 3390 1348 3394 1352
rect 3574 1348 3578 1352
rect 3638 1348 3642 1352
rect 3670 1348 3674 1352
rect 3702 1348 3706 1352
rect 3806 1348 3810 1352
rect 3822 1348 3826 1352
rect 3830 1348 3834 1352
rect 3878 1348 3882 1352
rect 3894 1348 3898 1352
rect 3926 1348 3930 1352
rect 3958 1348 3962 1352
rect 3998 1348 4002 1352
rect 54 1338 58 1342
rect 110 1338 114 1342
rect 246 1338 250 1342
rect 438 1338 442 1342
rect 574 1338 578 1342
rect 671 1338 675 1342
rect 702 1338 706 1342
rect 726 1338 730 1342
rect 742 1338 746 1342
rect 758 1338 762 1342
rect 846 1338 850 1342
rect 886 1338 890 1342
rect 934 1338 938 1342
rect 966 1338 970 1342
rect 1038 1338 1042 1342
rect 1054 1338 1058 1342
rect 1070 1338 1074 1342
rect 1094 1338 1098 1342
rect 1126 1338 1130 1342
rect 1142 1338 1146 1342
rect 1198 1338 1202 1342
rect 1230 1338 1234 1342
rect 1270 1338 1274 1342
rect 1302 1338 1306 1342
rect 1390 1338 1394 1342
rect 1454 1338 1458 1342
rect 1630 1338 1634 1342
rect 1686 1338 1690 1342
rect 1694 1338 1698 1342
rect 1742 1338 1746 1342
rect 1750 1338 1754 1342
rect 1814 1338 1818 1342
rect 1886 1338 1890 1342
rect 1894 1338 1898 1342
rect 1926 1338 1930 1342
rect 2214 1338 2218 1342
rect 2286 1338 2290 1342
rect 2318 1338 2322 1342
rect 2350 1338 2354 1342
rect 2374 1338 2378 1342
rect 2478 1338 2482 1342
rect 2486 1338 2490 1342
rect 2510 1338 2514 1342
rect 2526 1338 2530 1342
rect 2566 1338 2570 1342
rect 2654 1338 2658 1342
rect 2670 1338 2674 1342
rect 2718 1338 2722 1342
rect 2750 1338 2754 1342
rect 2774 1338 2778 1342
rect 2806 1338 2810 1342
rect 2838 1338 2842 1342
rect 2854 1338 2858 1342
rect 2886 1338 2890 1342
rect 2926 1338 2930 1342
rect 2942 1338 2946 1342
rect 2950 1338 2954 1342
rect 2990 1338 2994 1342
rect 3022 1338 3026 1342
rect 3166 1338 3170 1342
rect 3262 1338 3266 1342
rect 3278 1338 3282 1342
rect 3350 1338 3354 1342
rect 3358 1338 3362 1342
rect 3374 1338 3378 1342
rect 3398 1338 3402 1342
rect 3542 1338 3546 1342
rect 3630 1338 3634 1342
rect 3646 1338 3650 1342
rect 3694 1338 3698 1342
rect 3710 1338 3714 1342
rect 3734 1338 3738 1342
rect 3774 1338 3778 1342
rect 4038 1348 4042 1352
rect 4070 1348 4074 1352
rect 4102 1348 4106 1352
rect 4134 1348 4138 1352
rect 4166 1348 4170 1352
rect 4198 1348 4202 1352
rect 4214 1348 4218 1352
rect 4238 1348 4242 1352
rect 4262 1348 4266 1352
rect 4278 1348 4282 1352
rect 4302 1348 4306 1352
rect 4318 1348 4322 1352
rect 4350 1348 4354 1352
rect 3822 1338 3826 1342
rect 3870 1338 3874 1342
rect 4022 1338 4026 1342
rect 4094 1338 4098 1342
rect 4190 1338 4194 1342
rect 4254 1338 4258 1342
rect 4318 1338 4322 1342
rect 4374 1338 4378 1342
rect 230 1328 234 1332
rect 422 1328 426 1332
rect 590 1328 594 1332
rect 678 1328 682 1332
rect 1086 1328 1090 1332
rect 1334 1328 1338 1332
rect 1446 1328 1450 1332
rect 1566 1328 1570 1332
rect 1574 1328 1578 1332
rect 1638 1328 1642 1332
rect 1806 1328 1810 1332
rect 1846 1328 1850 1332
rect 1974 1328 1978 1332
rect 1990 1328 1994 1332
rect 2078 1328 2082 1332
rect 2198 1328 2202 1332
rect 2406 1328 2410 1332
rect 2526 1328 2530 1332
rect 2622 1328 2626 1332
rect 2646 1328 2650 1332
rect 2702 1328 2706 1332
rect 2758 1328 2762 1332
rect 2902 1328 2906 1332
rect 3150 1328 3154 1332
rect 3294 1328 3298 1332
rect 3422 1328 3426 1332
rect 3446 1328 3450 1332
rect 3526 1328 3530 1332
rect 3662 1328 3666 1332
rect 3750 1328 3754 1332
rect 3766 1328 3770 1332
rect 3854 1328 3858 1332
rect 4022 1328 4026 1332
rect 974 1318 978 1322
rect 1022 1318 1026 1322
rect 1102 1318 1106 1322
rect 1278 1318 1282 1322
rect 1310 1318 1314 1322
rect 1414 1318 1418 1322
rect 1478 1318 1482 1322
rect 1542 1318 1546 1322
rect 1606 1318 1610 1322
rect 1774 1318 1778 1322
rect 1854 1318 1858 1322
rect 2766 1318 2770 1322
rect 2790 1318 2794 1322
rect 3038 1318 3042 1322
rect 3070 1318 3074 1322
rect 3238 1318 3242 1322
rect 3614 1318 3618 1322
rect 3654 1318 3658 1322
rect 3726 1318 3730 1322
rect 3758 1318 3762 1322
rect 3790 1318 3794 1322
rect 4150 1318 4154 1322
rect 898 1303 902 1307
rect 905 1303 909 1307
rect 1930 1303 1934 1307
rect 1937 1303 1941 1307
rect 2954 1303 2958 1307
rect 2961 1303 2965 1307
rect 3978 1303 3982 1307
rect 3985 1303 3989 1307
rect 694 1288 698 1292
rect 750 1288 754 1292
rect 766 1288 770 1292
rect 838 1288 842 1292
rect 966 1288 970 1292
rect 1086 1288 1090 1292
rect 1150 1288 1154 1292
rect 1190 1288 1194 1292
rect 1358 1288 1362 1292
rect 1390 1288 1394 1292
rect 1710 1288 1714 1292
rect 1942 1288 1946 1292
rect 2070 1288 2074 1292
rect 2094 1288 2098 1292
rect 2718 1288 2722 1292
rect 2814 1288 2818 1292
rect 3142 1288 3146 1292
rect 3262 1288 3266 1292
rect 3454 1288 3458 1292
rect 3806 1288 3810 1292
rect 3862 1288 3866 1292
rect 3966 1288 3970 1292
rect 4094 1288 4098 1292
rect 4190 1288 4194 1292
rect 4286 1288 4290 1292
rect 4310 1288 4314 1292
rect 94 1278 98 1282
rect 262 1278 266 1282
rect 686 1278 690 1282
rect 758 1278 762 1282
rect 886 1278 890 1282
rect 1230 1278 1234 1282
rect 1350 1278 1354 1282
rect 1438 1278 1442 1282
rect 1606 1278 1610 1282
rect 110 1268 114 1272
rect 246 1268 250 1272
rect 358 1268 362 1272
rect 374 1268 378 1272
rect 390 1268 394 1272
rect 430 1268 434 1272
rect 582 1268 586 1272
rect 614 1268 618 1272
rect 638 1268 642 1272
rect 662 1268 666 1272
rect 710 1268 714 1272
rect 734 1268 738 1272
rect 742 1268 746 1272
rect 790 1268 794 1272
rect 854 1268 858 1272
rect 870 1268 874 1272
rect 910 1268 914 1272
rect 926 1268 930 1272
rect 942 1268 946 1272
rect 950 1268 954 1272
rect 974 1268 978 1272
rect 1094 1268 1098 1272
rect 1102 1268 1106 1272
rect 1126 1268 1130 1272
rect 1158 1268 1162 1272
rect 1182 1268 1186 1272
rect 1214 1268 1218 1272
rect 1262 1268 1266 1272
rect 1286 1268 1290 1272
rect 1318 1268 1322 1272
rect 1366 1268 1370 1272
rect 1398 1268 1402 1272
rect 1446 1268 1450 1272
rect 1502 1268 1506 1272
rect 1534 1268 1538 1272
rect 1542 1268 1546 1272
rect 1574 1268 1578 1272
rect 1622 1268 1626 1272
rect 1646 1268 1650 1272
rect 1766 1278 1770 1282
rect 1774 1278 1778 1282
rect 1878 1278 1882 1282
rect 2014 1278 2018 1282
rect 2062 1278 2066 1282
rect 2190 1278 2194 1282
rect 2406 1278 2410 1282
rect 2518 1278 2522 1282
rect 2614 1278 2618 1282
rect 2774 1278 2778 1282
rect 2830 1278 2834 1282
rect 2910 1278 2914 1282
rect 3070 1278 3074 1282
rect 1702 1268 1706 1272
rect 1718 1268 1722 1272
rect 1782 1268 1786 1272
rect 1902 1268 1906 1272
rect 1934 1268 1938 1272
rect 2022 1268 2026 1272
rect 2054 1268 2058 1272
rect 2078 1268 2082 1272
rect 2206 1268 2210 1272
rect 2278 1268 2282 1272
rect 2294 1268 2298 1272
rect 2422 1268 2426 1272
rect 2510 1268 2514 1272
rect 2630 1268 2634 1272
rect 2710 1268 2714 1272
rect 2726 1268 2730 1272
rect 2742 1268 2746 1272
rect 2790 1268 2794 1272
rect 2806 1268 2810 1272
rect 2926 1268 2930 1272
rect 3014 1268 3018 1272
rect 3046 1268 3050 1272
rect 3086 1268 3090 1272
rect 3134 1268 3138 1272
rect 3174 1268 3178 1272
rect 3246 1268 3250 1272
rect 3254 1268 3258 1272
rect 3302 1278 3306 1282
rect 3374 1278 3378 1282
rect 3422 1278 3426 1282
rect 3286 1268 3290 1272
rect 3302 1268 3306 1272
rect 3318 1268 3322 1272
rect 3358 1268 3362 1272
rect 3382 1268 3386 1272
rect 3398 1268 3402 1272
rect 3414 1268 3418 1272
rect 3446 1268 3450 1272
rect 3462 1268 3466 1272
rect 3470 1268 3474 1272
rect 3534 1268 3538 1272
rect 3646 1278 3650 1282
rect 3686 1278 3690 1282
rect 3726 1278 3730 1282
rect 3774 1278 3778 1282
rect 3814 1278 3818 1282
rect 3878 1278 3882 1282
rect 3926 1278 3930 1282
rect 4022 1278 4026 1282
rect 4102 1278 4106 1282
rect 4198 1278 4202 1282
rect 4254 1278 4258 1282
rect 4294 1278 4298 1282
rect 3614 1268 3618 1272
rect 3694 1268 3698 1272
rect 3742 1268 3746 1272
rect 3782 1268 3786 1272
rect 3830 1268 3834 1272
rect 4086 1268 4090 1272
rect 4278 1268 4282 1272
rect 4318 1268 4322 1272
rect 158 1258 162 1262
rect 198 1258 202 1262
rect 446 1258 450 1262
rect 462 1258 466 1262
rect 494 1258 498 1262
rect 526 1258 530 1262
rect 558 1258 562 1262
rect 590 1258 594 1262
rect 606 1258 610 1262
rect 630 1258 634 1262
rect 670 1258 674 1262
rect 782 1258 786 1262
rect 798 1258 802 1262
rect 822 1258 826 1262
rect 830 1258 834 1262
rect 862 1258 866 1262
rect 878 1258 882 1262
rect 918 1258 922 1262
rect 934 1258 938 1262
rect 1046 1258 1050 1262
rect 1134 1258 1138 1262
rect 1190 1258 1194 1262
rect 1206 1258 1210 1262
rect 1246 1258 1250 1262
rect 1278 1258 1282 1262
rect 1294 1258 1298 1262
rect 1326 1258 1330 1262
rect 1374 1258 1378 1262
rect 1406 1258 1410 1262
rect 1462 1258 1466 1262
rect 1478 1258 1482 1262
rect 1502 1258 1506 1262
rect 1510 1258 1514 1262
rect 1526 1258 1530 1262
rect 1550 1258 1554 1262
rect 1566 1258 1570 1262
rect 1582 1258 1586 1262
rect 1630 1258 1634 1262
rect 1638 1258 1642 1262
rect 1654 1258 1658 1262
rect 1670 1258 1674 1262
rect 1694 1258 1698 1262
rect 1734 1258 1738 1262
rect 1758 1258 1762 1262
rect 1790 1258 1794 1262
rect 1814 1258 1818 1262
rect 1822 1258 1826 1262
rect 1838 1258 1842 1262
rect 1862 1258 1866 1262
rect 1894 1258 1898 1262
rect 1910 1258 1914 1262
rect 1950 1258 1954 1262
rect 1982 1258 1986 1262
rect 1990 1258 1994 1262
rect 1998 1258 2002 1262
rect 2014 1258 2018 1262
rect 2062 1258 2066 1262
rect 2150 1258 2154 1262
rect 2294 1258 2298 1262
rect 2462 1258 2466 1262
rect 2478 1258 2482 1262
rect 2533 1258 2537 1262
rect 2670 1258 2674 1262
rect 2678 1258 2682 1262
rect 2702 1258 2706 1262
rect 2742 1258 2746 1262
rect 2750 1258 2754 1262
rect 2798 1258 2802 1262
rect 2870 1258 2874 1262
rect 3038 1258 3042 1262
rect 3054 1258 3058 1262
rect 3094 1258 3098 1262
rect 3102 1258 3106 1262
rect 3174 1258 3178 1262
rect 3182 1258 3186 1262
rect 3230 1258 3234 1262
rect 3238 1258 3242 1262
rect 3278 1258 3282 1262
rect 3310 1258 3314 1262
rect 3326 1258 3330 1262
rect 3350 1258 3354 1262
rect 3406 1258 3410 1262
rect 3438 1258 3442 1262
rect 3478 1258 3482 1262
rect 3502 1258 3506 1262
rect 3518 1258 3522 1262
rect 3526 1258 3530 1262
rect 3542 1258 3546 1262
rect 3582 1258 3586 1262
rect 3606 1258 3610 1262
rect 3622 1258 3626 1262
rect 3670 1258 3674 1262
rect 3702 1258 3706 1262
rect 3750 1258 3754 1262
rect 3758 1258 3762 1262
rect 3790 1258 3794 1262
rect 3838 1258 3842 1262
rect 3846 1258 3850 1262
rect 3894 1258 3898 1262
rect 3910 1258 3914 1262
rect 3942 1258 3946 1262
rect 3998 1258 4002 1262
rect 4022 1258 4026 1262
rect 4054 1258 4058 1262
rect 4110 1258 4114 1262
rect 4150 1258 4154 1262
rect 4174 1258 4178 1262
rect 4214 1258 4218 1262
rect 4230 1258 4234 1262
rect 4254 1258 4258 1262
rect 4270 1258 4274 1262
rect 4326 1258 4330 1262
rect 4342 1258 4346 1262
rect 4366 1258 4370 1262
rect 142 1250 146 1254
rect 198 1248 202 1252
rect 414 1248 418 1252
rect 454 1248 458 1252
rect 486 1248 490 1252
rect 518 1248 522 1252
rect 550 1248 554 1252
rect 614 1248 618 1252
rect 646 1248 650 1252
rect 838 1248 842 1252
rect 1078 1248 1082 1252
rect 1118 1248 1122 1252
rect 1150 1248 1154 1252
rect 1174 1248 1178 1252
rect 1310 1248 1314 1252
rect 1342 1248 1346 1252
rect 1390 1248 1394 1252
rect 1422 1248 1426 1252
rect 1494 1248 1498 1252
rect 1510 1248 1514 1252
rect 1566 1248 1570 1252
rect 1598 1248 1602 1252
rect 1934 1248 1938 1252
rect 2094 1248 2098 1252
rect 2238 1250 2242 1254
rect 2470 1248 2474 1252
rect 2662 1250 2666 1254
rect 2750 1248 2754 1252
rect 2974 1248 2978 1252
rect 3110 1248 3114 1252
rect 3126 1248 3130 1252
rect 3150 1248 3154 1252
rect 3166 1248 3170 1252
rect 3214 1248 3218 1252
rect 3326 1248 3330 1252
rect 3342 1248 3346 1252
rect 3374 1248 3378 1252
rect 3902 1248 3906 1252
rect 3934 1248 3938 1252
rect 4006 1248 4010 1252
rect 4014 1248 4018 1252
rect 4046 1248 4050 1252
rect 4126 1248 4130 1252
rect 4142 1248 4146 1252
rect 4206 1248 4210 1252
rect 4262 1248 4266 1252
rect 4334 1248 4338 1252
rect 4358 1248 4362 1252
rect 470 1238 474 1242
rect 502 1238 506 1242
rect 534 1238 538 1242
rect 566 1238 570 1242
rect 662 1238 666 1242
rect 694 1238 698 1242
rect 710 1238 714 1242
rect 734 1238 738 1242
rect 966 1238 970 1242
rect 1158 1238 1162 1242
rect 1622 1238 1626 1242
rect 2110 1238 2114 1242
rect 3382 1238 3386 1242
rect 3918 1238 3922 1242
rect 3950 1238 3954 1242
rect 3990 1238 3994 1242
rect 4030 1238 4034 1242
rect 4062 1238 4066 1242
rect 4158 1238 4162 1242
rect 4222 1238 4226 1242
rect 4246 1238 4250 1242
rect 4350 1238 4354 1242
rect 366 1228 370 1232
rect 1846 1228 1850 1232
rect 2326 1228 2330 1232
rect 2662 1227 2666 1231
rect 3230 1228 3234 1232
rect 3502 1228 3506 1232
rect 14 1218 18 1222
rect 142 1218 146 1222
rect 198 1218 202 1222
rect 462 1218 466 1222
rect 494 1218 498 1222
rect 526 1218 530 1222
rect 558 1218 562 1222
rect 654 1218 658 1222
rect 750 1218 754 1222
rect 814 1218 818 1222
rect 1030 1218 1034 1222
rect 1062 1218 1066 1222
rect 1110 1218 1114 1222
rect 1294 1218 1298 1222
rect 1326 1218 1330 1222
rect 1582 1218 1586 1222
rect 1742 1218 1746 1222
rect 2238 1218 2242 1222
rect 2302 1218 2306 1222
rect 2470 1218 2474 1222
rect 2974 1218 2978 1222
rect 3022 1218 3026 1222
rect 3198 1218 3202 1222
rect 3566 1218 3570 1222
rect 3590 1218 3594 1222
rect 3622 1218 3626 1222
rect 3654 1218 3658 1222
rect 3670 1218 3674 1222
rect 3702 1218 3706 1222
rect 3766 1218 3770 1222
rect 3862 1218 3866 1222
rect 3894 1218 3898 1222
rect 3998 1218 4002 1222
rect 4382 1218 4386 1222
rect 394 1203 398 1207
rect 401 1203 405 1207
rect 1418 1203 1422 1207
rect 1425 1203 1429 1207
rect 2442 1203 2446 1207
rect 2449 1203 2453 1207
rect 3474 1203 3478 1207
rect 3481 1203 3485 1207
rect 38 1188 42 1192
rect 110 1188 114 1192
rect 206 1188 210 1192
rect 614 1188 618 1192
rect 790 1188 794 1192
rect 942 1188 946 1192
rect 1310 1188 1314 1192
rect 1358 1188 1362 1192
rect 1502 1188 1506 1192
rect 1518 1188 1522 1192
rect 1550 1188 1554 1192
rect 1614 1188 1618 1192
rect 1678 1188 1682 1192
rect 1798 1188 1802 1192
rect 1910 1188 1914 1192
rect 2190 1188 2194 1192
rect 2494 1188 2498 1192
rect 3126 1188 3130 1192
rect 3278 1188 3282 1192
rect 3374 1188 3378 1192
rect 3438 1188 3442 1192
rect 3510 1188 3514 1192
rect 3670 1188 3674 1192
rect 3990 1188 3994 1192
rect 4022 1188 4026 1192
rect 4110 1188 4114 1192
rect 4134 1188 4138 1192
rect 4166 1188 4170 1192
rect 4246 1188 4250 1192
rect 4270 1188 4274 1192
rect 4310 1188 4314 1192
rect 4358 1188 4362 1192
rect 398 1178 402 1182
rect 582 1178 586 1182
rect 1182 1179 1186 1183
rect 2150 1179 2154 1183
rect 2622 1178 2626 1182
rect 2766 1179 2770 1183
rect 3214 1178 3218 1182
rect 4214 1178 4218 1182
rect 350 1168 354 1172
rect 574 1168 578 1172
rect 646 1168 650 1172
rect 870 1168 874 1172
rect 918 1168 922 1172
rect 926 1168 930 1172
rect 1438 1168 1442 1172
rect 3966 1168 3970 1172
rect 4014 1168 4018 1172
rect 4046 1168 4050 1172
rect 4102 1168 4106 1172
rect 4174 1168 4178 1172
rect 4206 1168 4210 1172
rect 4238 1168 4242 1172
rect 4262 1168 4266 1172
rect 4302 1168 4306 1172
rect 4326 1168 4330 1172
rect 4334 1168 4338 1172
rect 4366 1168 4370 1172
rect 150 1158 154 1162
rect 206 1158 210 1162
rect 422 1158 426 1162
rect 430 1158 434 1162
rect 486 1158 490 1162
rect 518 1158 522 1162
rect 550 1158 554 1162
rect 566 1158 570 1162
rect 574 1158 578 1162
rect 662 1158 666 1162
rect 694 1158 698 1162
rect 838 1158 842 1162
rect 862 1158 866 1162
rect 1102 1158 1106 1162
rect 1182 1156 1186 1160
rect 1350 1158 1354 1162
rect 1566 1158 1570 1162
rect 1630 1158 1634 1162
rect 1662 1158 1666 1162
rect 1726 1158 1730 1162
rect 1734 1158 1738 1162
rect 1846 1158 1850 1162
rect 1886 1158 1890 1162
rect 1974 1158 1978 1162
rect 1990 1158 1994 1162
rect 2150 1156 2154 1160
rect 2238 1158 2242 1162
rect 2270 1158 2274 1162
rect 2494 1158 2498 1162
rect 2574 1158 2578 1162
rect 2766 1156 2770 1160
rect 2838 1158 2842 1162
rect 2870 1158 2874 1162
rect 2902 1158 2906 1162
rect 2934 1158 2938 1162
rect 3022 1158 3026 1162
rect 3038 1158 3042 1162
rect 3054 1158 3058 1162
rect 3086 1158 3090 1162
rect 3174 1158 3178 1162
rect 3478 1158 3482 1162
rect 3670 1158 3674 1162
rect 3710 1158 3714 1162
rect 3806 1158 3810 1162
rect 3950 1158 3954 1162
rect 3998 1158 4002 1162
rect 4030 1158 4034 1162
rect 4054 1158 4058 1162
rect 4118 1158 4122 1162
rect 4150 1158 4154 1162
rect 4158 1158 4162 1162
rect 4190 1158 4194 1162
rect 4222 1158 4226 1162
rect 4294 1158 4298 1162
rect 4318 1158 4322 1162
rect 4350 1158 4354 1162
rect 22 1148 26 1152
rect 86 1148 90 1152
rect 94 1148 98 1152
rect 126 1148 130 1152
rect 142 1148 146 1152
rect 182 1148 186 1152
rect 206 1148 210 1152
rect 310 1148 314 1152
rect 382 1148 386 1152
rect 446 1148 450 1152
rect 454 1148 458 1152
rect 502 1148 506 1152
rect 534 1148 538 1152
rect 582 1148 586 1152
rect 630 1148 634 1152
rect 646 1148 650 1152
rect 678 1148 682 1152
rect 710 1148 714 1152
rect 726 1148 730 1152
rect 750 1148 754 1152
rect 766 1148 770 1152
rect 806 1148 810 1152
rect 822 1148 826 1152
rect 918 1148 922 1152
rect 958 1148 962 1152
rect 982 1148 986 1152
rect 1006 1148 1010 1152
rect 1038 1148 1042 1152
rect 1054 1148 1058 1152
rect 1070 1148 1074 1152
rect 1118 1148 1122 1152
rect 1142 1148 1146 1152
rect 1166 1148 1170 1152
rect 1334 1148 1338 1152
rect 1422 1148 1426 1152
rect 1454 1148 1458 1152
rect 1494 1148 1498 1152
rect 1518 1148 1522 1152
rect 1550 1148 1554 1152
rect 1574 1148 1578 1152
rect 1614 1148 1618 1152
rect 1646 1148 1650 1152
rect 1670 1148 1674 1152
rect 1702 1148 1706 1152
rect 1710 1148 1714 1152
rect 1758 1148 1762 1152
rect 1814 1148 1818 1152
rect 1830 1148 1834 1152
rect 1854 1148 1858 1152
rect 1878 1148 1882 1152
rect 1902 1148 1906 1152
rect 1966 1148 1970 1152
rect 1974 1148 1978 1152
rect 1998 1148 2002 1152
rect 2166 1148 2170 1152
rect 2190 1148 2194 1152
rect 2222 1148 2226 1152
rect 2254 1148 2258 1152
rect 2262 1148 2266 1152
rect 2278 1148 2282 1152
rect 2310 1148 2314 1152
rect 2390 1148 2394 1152
rect 2478 1148 2482 1152
rect 2558 1148 2562 1152
rect 2582 1148 2586 1152
rect 2637 1148 2641 1152
rect 2678 1148 2682 1152
rect 2806 1148 2810 1152
rect 2838 1148 2842 1152
rect 2854 1148 2858 1152
rect 2878 1148 2882 1152
rect 2918 1148 2922 1152
rect 2950 1148 2954 1152
rect 2990 1148 2994 1152
rect 3006 1148 3010 1152
rect 3070 1148 3074 1152
rect 3102 1148 3106 1152
rect 3134 1148 3138 1152
rect 3142 1148 3146 1152
rect 3190 1148 3194 1152
rect 3222 1148 3226 1152
rect 3254 1148 3258 1152
rect 3286 1148 3290 1152
rect 3294 1148 3298 1152
rect 3318 1148 3322 1152
rect 3326 1148 3330 1152
rect 3358 1148 3362 1152
rect 3374 1148 3378 1152
rect 3422 1148 3426 1152
rect 3454 1148 3458 1152
rect 3670 1148 3674 1152
rect 3726 1148 3730 1152
rect 3742 1148 3746 1152
rect 3782 1148 3786 1152
rect 3822 1148 3826 1152
rect 3846 1148 3850 1152
rect 3926 1148 3930 1152
rect 3958 1148 3962 1152
rect 4006 1148 4010 1152
rect 4038 1148 4042 1152
rect 4062 1148 4066 1152
rect 4110 1148 4114 1152
rect 4134 1148 4138 1152
rect 4166 1148 4170 1152
rect 4198 1148 4202 1152
rect 4230 1148 4234 1152
rect 4270 1148 4274 1152
rect 4294 1148 4298 1152
rect 4326 1148 4330 1152
rect 4358 1148 4362 1152
rect 62 1138 66 1142
rect 126 1138 130 1142
rect 158 1138 162 1142
rect 254 1138 258 1142
rect 366 1138 370 1142
rect 382 1138 386 1142
rect 414 1138 418 1142
rect 462 1138 466 1142
rect 478 1138 482 1142
rect 494 1138 498 1142
rect 526 1138 530 1142
rect 558 1138 562 1142
rect 606 1138 610 1142
rect 638 1138 642 1142
rect 670 1138 674 1142
rect 686 1138 690 1142
rect 702 1138 706 1142
rect 742 1138 746 1142
rect 774 1138 778 1142
rect 814 1138 818 1142
rect 846 1138 850 1142
rect 902 1138 906 1142
rect 958 1138 962 1142
rect 990 1138 994 1142
rect 1046 1138 1050 1142
rect 1078 1138 1082 1142
rect 1086 1138 1090 1142
rect 1102 1138 1106 1142
rect 1110 1138 1114 1142
rect 1142 1138 1146 1142
rect 1214 1138 1218 1142
rect 1318 1138 1322 1142
rect 1454 1138 1458 1142
rect 1478 1138 1482 1142
rect 1542 1138 1546 1142
rect 1606 1138 1610 1142
rect 1638 1138 1642 1142
rect 1694 1138 1698 1142
rect 1790 1138 1794 1142
rect 1822 1138 1826 1142
rect 1870 1138 1874 1142
rect 1958 1138 1962 1142
rect 1998 1138 2002 1142
rect 2014 1138 2018 1142
rect 2118 1138 2122 1142
rect 2214 1138 2218 1142
rect 2246 1138 2250 1142
rect 2286 1138 2290 1142
rect 2318 1138 2322 1142
rect 2446 1138 2450 1142
rect 2534 1138 2538 1142
rect 2550 1138 2554 1142
rect 2614 1138 2618 1142
rect 2734 1138 2738 1142
rect 2830 1138 2834 1142
rect 2862 1138 2866 1142
rect 2894 1138 2898 1142
rect 2926 1138 2930 1142
rect 2974 1138 2978 1142
rect 2982 1138 2986 1142
rect 3014 1138 3018 1142
rect 3046 1138 3050 1142
rect 3078 1138 3082 1142
rect 3094 1138 3098 1142
rect 3110 1138 3114 1142
rect 3134 1138 3138 1142
rect 3150 1138 3154 1142
rect 3198 1138 3202 1142
rect 3206 1138 3210 1142
rect 3230 1138 3234 1142
rect 3254 1138 3258 1142
rect 3262 1138 3266 1142
rect 3278 1138 3282 1142
rect 3302 1138 3306 1142
rect 3334 1138 3338 1142
rect 3350 1138 3354 1142
rect 3366 1138 3370 1142
rect 3414 1138 3418 1142
rect 3494 1138 3498 1142
rect 3502 1138 3506 1142
rect 3622 1138 3626 1142
rect 3734 1138 3738 1142
rect 3774 1138 3778 1142
rect 3790 1138 3794 1142
rect 3798 1138 3802 1142
rect 3814 1138 3818 1142
rect 3830 1138 3834 1142
rect 3838 1138 3842 1142
rect 3886 1138 3890 1142
rect 4070 1138 4074 1142
rect 4086 1138 4090 1142
rect 4126 1138 4130 1142
rect 270 1128 274 1132
rect 950 1128 954 1132
rect 1006 1128 1010 1132
rect 1230 1128 1234 1132
rect 1366 1128 1370 1132
rect 1494 1128 1498 1132
rect 1534 1128 1538 1132
rect 1590 1128 1594 1132
rect 1670 1128 1674 1132
rect 1726 1128 1730 1132
rect 1742 1128 1746 1132
rect 1870 1128 1874 1132
rect 1894 1128 1898 1132
rect 1918 1128 1922 1132
rect 1942 1128 1946 1132
rect 2102 1128 2106 1132
rect 2206 1128 2210 1132
rect 2238 1128 2242 1132
rect 2302 1128 2306 1132
rect 2334 1128 2338 1132
rect 2430 1128 2434 1132
rect 2606 1128 2610 1132
rect 2718 1128 2722 1132
rect 2822 1128 2826 1132
rect 3118 1128 3122 1132
rect 3238 1128 3242 1132
rect 3398 1128 3402 1132
rect 3470 1128 3474 1132
rect 3606 1128 3610 1132
rect 3702 1128 3706 1132
rect 3742 1128 3746 1132
rect 3758 1128 3762 1132
rect 3870 1128 3874 1132
rect 3902 1128 3906 1132
rect 3942 1128 3946 1132
rect 4086 1128 4090 1132
rect 430 1118 434 1122
rect 518 1118 522 1122
rect 550 1118 554 1122
rect 710 1118 714 1122
rect 766 1118 770 1122
rect 838 1118 842 1122
rect 862 1118 866 1122
rect 982 1118 986 1122
rect 1022 1118 1026 1122
rect 1070 1118 1074 1122
rect 1118 1118 1122 1122
rect 1350 1118 1354 1122
rect 1382 1118 1386 1122
rect 1470 1118 1474 1122
rect 1750 1118 1754 1122
rect 1846 1118 1850 1122
rect 1950 1118 1954 1122
rect 2022 1118 2026 1122
rect 2294 1118 2298 1122
rect 2326 1118 2330 1122
rect 2350 1118 2354 1122
rect 2542 1118 2546 1122
rect 2598 1118 2602 1122
rect 2814 1118 2818 1122
rect 2934 1118 2938 1122
rect 3006 1118 3010 1122
rect 3158 1118 3162 1122
rect 3342 1118 3346 1122
rect 3526 1118 3530 1122
rect 3694 1118 3698 1122
rect 3710 1118 3714 1122
rect 3766 1118 3770 1122
rect 3862 1118 3866 1122
rect 3878 1118 3882 1122
rect 898 1103 902 1107
rect 905 1103 909 1107
rect 1930 1103 1934 1107
rect 1937 1103 1941 1107
rect 2954 1103 2958 1107
rect 2961 1103 2965 1107
rect 3978 1103 3982 1107
rect 3985 1103 3989 1107
rect 270 1088 274 1092
rect 614 1088 618 1092
rect 934 1088 938 1092
rect 998 1088 1002 1092
rect 1254 1088 1258 1092
rect 1358 1088 1362 1092
rect 1398 1088 1402 1092
rect 1566 1088 1570 1092
rect 1622 1088 1626 1092
rect 1734 1088 1738 1092
rect 2022 1088 2026 1092
rect 2062 1088 2066 1092
rect 2390 1088 2394 1092
rect 2462 1088 2466 1092
rect 2558 1088 2562 1092
rect 2574 1088 2578 1092
rect 2614 1088 2618 1092
rect 2894 1088 2898 1092
rect 3246 1088 3250 1092
rect 3286 1088 3290 1092
rect 3350 1088 3354 1092
rect 3462 1088 3466 1092
rect 3558 1088 3562 1092
rect 3718 1088 3722 1092
rect 3734 1088 3738 1092
rect 4094 1088 4098 1092
rect 4118 1088 4122 1092
rect 4254 1088 4258 1092
rect 4262 1088 4266 1092
rect 4302 1088 4306 1092
rect 4342 1088 4346 1092
rect 4374 1088 4378 1092
rect 6 1078 10 1082
rect 142 1078 146 1082
rect 350 1078 354 1082
rect 534 1078 538 1082
rect 854 1078 858 1082
rect 966 1078 970 1082
rect 982 1078 986 1082
rect 1174 1078 1178 1082
rect 1390 1078 1394 1082
rect 1422 1078 1426 1082
rect 1534 1078 1538 1082
rect 1758 1078 1762 1082
rect 1806 1078 1810 1082
rect 1854 1078 1858 1082
rect 1902 1078 1906 1082
rect 1974 1078 1978 1082
rect 2030 1078 2034 1082
rect 2134 1078 2138 1082
rect 2174 1078 2178 1082
rect 2262 1078 2266 1082
rect 2382 1078 2386 1082
rect 2422 1078 2426 1082
rect 2534 1078 2538 1082
rect 2758 1078 2762 1082
rect 2846 1078 2850 1082
rect 2886 1078 2890 1082
rect 2966 1078 2970 1082
rect 3094 1078 3098 1082
rect 3206 1078 3210 1082
rect 3254 1078 3258 1082
rect 3398 1078 3402 1082
rect 3478 1078 3482 1082
rect 3574 1078 3578 1082
rect 3630 1078 3634 1082
rect 3662 1078 3666 1082
rect 3702 1078 3706 1082
rect 3838 1078 3842 1082
rect 3974 1078 3978 1082
rect 4126 1078 4130 1082
rect 4150 1078 4154 1082
rect 4190 1078 4194 1082
rect 4206 1078 4210 1082
rect 30 1068 34 1072
rect 158 1068 162 1072
rect 230 1068 234 1072
rect 366 1068 370 1072
rect 518 1068 522 1072
rect 646 1068 650 1072
rect 742 1068 746 1072
rect 838 1068 842 1072
rect 1006 1068 1010 1072
rect 1022 1068 1026 1072
rect 1046 1068 1050 1072
rect 1158 1068 1162 1072
rect 1310 1068 1314 1072
rect 1350 1068 1354 1072
rect 1374 1068 1378 1072
rect 1382 1068 1386 1072
rect 1470 1068 1474 1072
rect 22 1058 26 1062
rect 198 1058 202 1062
rect 230 1058 234 1062
rect 254 1058 258 1062
rect 310 1058 314 1062
rect 470 1058 474 1062
rect 654 1058 658 1062
rect 686 1058 690 1062
rect 718 1058 722 1062
rect 750 1058 754 1062
rect 894 1058 898 1062
rect 982 1058 986 1062
rect 1014 1058 1018 1062
rect 1022 1058 1026 1062
rect 1054 1058 1058 1062
rect 1070 1058 1074 1062
rect 1102 1058 1106 1062
rect 1110 1058 1114 1062
rect 1270 1058 1274 1062
rect 1278 1058 1282 1062
rect 1302 1058 1306 1062
rect 1326 1058 1330 1062
rect 1334 1058 1338 1062
rect 1342 1058 1346 1062
rect 1430 1058 1434 1062
rect 1438 1058 1442 1062
rect 1462 1058 1466 1062
rect 1470 1058 1474 1062
rect 1542 1068 1546 1072
rect 1574 1068 1578 1072
rect 1606 1068 1610 1072
rect 1630 1068 1634 1072
rect 1646 1068 1650 1072
rect 1686 1068 1690 1072
rect 1694 1068 1698 1072
rect 1710 1068 1714 1072
rect 1782 1068 1786 1072
rect 1814 1068 1818 1072
rect 1822 1068 1826 1072
rect 1838 1068 1842 1072
rect 1878 1068 1882 1072
rect 1910 1068 1914 1072
rect 1934 1068 1938 1072
rect 1990 1068 1994 1072
rect 2094 1068 2098 1072
rect 2110 1068 2114 1072
rect 2134 1068 2138 1072
rect 2278 1068 2282 1072
rect 2350 1068 2354 1072
rect 2478 1068 2482 1072
rect 2550 1068 2554 1072
rect 2638 1068 2642 1072
rect 2654 1068 2658 1072
rect 2677 1068 2681 1072
rect 2774 1068 2778 1072
rect 2918 1068 2922 1072
rect 2950 1068 2954 1072
rect 2990 1068 2994 1072
rect 3110 1068 3114 1072
rect 3198 1068 3202 1072
rect 3222 1068 3226 1072
rect 3238 1068 3242 1072
rect 3262 1068 3266 1072
rect 3302 1068 3306 1072
rect 3326 1068 3330 1072
rect 3358 1068 3362 1072
rect 3406 1068 3410 1072
rect 3438 1068 3442 1072
rect 3510 1068 3514 1072
rect 3518 1068 3522 1072
rect 3542 1068 3546 1072
rect 3558 1068 3562 1072
rect 3566 1068 3570 1072
rect 3622 1068 3626 1072
rect 3646 1068 3650 1072
rect 3662 1068 3666 1072
rect 3726 1068 3730 1072
rect 3742 1068 3746 1072
rect 3854 1068 3858 1072
rect 3950 1068 3954 1072
rect 4110 1068 4114 1072
rect 4174 1068 4178 1072
rect 4294 1068 4298 1072
rect 1486 1058 1490 1062
rect 1502 1058 1506 1062
rect 1518 1058 1522 1062
rect 1534 1058 1538 1062
rect 1582 1058 1586 1062
rect 1638 1058 1642 1062
rect 1654 1058 1658 1062
rect 1670 1058 1674 1062
rect 1702 1058 1706 1062
rect 1750 1058 1754 1062
rect 1774 1058 1778 1062
rect 1782 1058 1786 1062
rect 1806 1058 1810 1062
rect 1830 1058 1834 1062
rect 1870 1058 1874 1062
rect 1878 1058 1882 1062
rect 1902 1058 1906 1062
rect 1942 1058 1946 1062
rect 1958 1058 1962 1062
rect 1990 1058 1994 1062
rect 2006 1058 2010 1062
rect 2046 1058 2050 1062
rect 2118 1058 2122 1062
rect 2142 1058 2146 1062
rect 2150 1058 2154 1062
rect 2222 1058 2226 1062
rect 2318 1058 2322 1062
rect 2358 1058 2362 1062
rect 2366 1058 2370 1062
rect 2398 1058 2402 1062
rect 2430 1058 2434 1062
rect 2438 1058 2442 1062
rect 2598 1058 2602 1062
rect 2630 1058 2634 1062
rect 2662 1058 2666 1062
rect 2718 1058 2722 1062
rect 2862 1058 2866 1062
rect 2870 1058 2874 1062
rect 2886 1058 2890 1062
rect 2942 1058 2946 1062
rect 2998 1058 3002 1062
rect 3110 1058 3114 1062
rect 3182 1058 3186 1062
rect 3206 1058 3210 1062
rect 3222 1058 3226 1062
rect 3270 1058 3274 1062
rect 3334 1058 3338 1062
rect 3366 1058 3370 1062
rect 3430 1058 3434 1062
rect 3446 1058 3450 1062
rect 3502 1058 3506 1062
rect 3534 1058 3538 1062
rect 3566 1058 3570 1062
rect 3598 1058 3602 1062
rect 3670 1058 3674 1062
rect 3686 1058 3690 1062
rect 3798 1058 3802 1062
rect 3934 1058 3938 1062
rect 3974 1058 3978 1062
rect 4014 1058 4018 1062
rect 4046 1058 4050 1062
rect 4078 1058 4082 1062
rect 4102 1058 4106 1062
rect 4150 1058 4154 1062
rect 4166 1058 4170 1062
rect 4190 1058 4194 1062
rect 4206 1058 4210 1062
rect 4238 1058 4242 1062
rect 4278 1058 4282 1062
rect 4318 1058 4322 1062
rect 4326 1058 4330 1062
rect 4358 1058 4362 1062
rect 206 1048 210 1052
rect 414 1048 418 1052
rect 422 1048 426 1052
rect 486 1050 490 1054
rect 654 1048 658 1052
rect 670 1048 674 1052
rect 678 1048 682 1052
rect 710 1048 714 1052
rect 750 1048 754 1052
rect 766 1048 770 1052
rect 790 1048 794 1052
rect 1062 1048 1066 1052
rect 1110 1048 1114 1052
rect 1358 1048 1362 1052
rect 1502 1048 1506 1052
rect 1566 1048 1570 1052
rect 1582 1048 1586 1052
rect 1598 1048 1602 1052
rect 1622 1048 1626 1052
rect 1654 1048 1658 1052
rect 1718 1048 1722 1052
rect 1846 1048 1850 1052
rect 2022 1048 2026 1052
rect 2078 1048 2082 1052
rect 2310 1050 2314 1054
rect 2374 1048 2378 1052
rect 2654 1048 2658 1052
rect 2806 1050 2810 1054
rect 2894 1048 2898 1052
rect 2926 1048 2930 1052
rect 2966 1048 2970 1052
rect 3142 1050 3146 1054
rect 3286 1048 3290 1052
rect 3294 1048 3298 1052
rect 3350 1048 3354 1052
rect 3366 1048 3370 1052
rect 3382 1048 3386 1052
rect 3462 1048 3466 1052
rect 3486 1048 3490 1052
rect 3606 1048 3610 1052
rect 3710 1048 3714 1052
rect 3886 1050 3890 1054
rect 3926 1048 3930 1052
rect 3982 1048 3986 1052
rect 4006 1048 4010 1052
rect 4038 1048 4042 1052
rect 4070 1048 4074 1052
rect 4158 1048 4162 1052
rect 4198 1048 4202 1052
rect 4230 1048 4234 1052
rect 4262 1048 4266 1052
rect 694 1038 698 1042
rect 726 1038 730 1042
rect 1078 1038 1082 1042
rect 1774 1038 1778 1042
rect 1870 1038 1874 1042
rect 3942 1038 3946 1042
rect 3966 1038 3970 1042
rect 3974 1038 3978 1042
rect 4022 1038 4026 1042
rect 4054 1038 4058 1042
rect 4086 1038 4090 1042
rect 4142 1038 4146 1042
rect 4214 1038 4218 1042
rect 4246 1038 4250 1042
rect 486 1027 490 1031
rect 1046 1028 1050 1032
rect 2310 1027 2314 1031
rect 2806 1027 2810 1031
rect 3014 1028 3018 1032
rect 3142 1027 3146 1031
rect 3886 1027 3890 1031
rect 206 1018 210 1022
rect 414 1018 418 1022
rect 686 1018 690 1022
rect 718 1018 722 1022
rect 790 1018 794 1022
rect 982 1018 986 1022
rect 1086 1018 1090 1022
rect 1110 1018 1114 1022
rect 1294 1018 1298 1022
rect 1958 1018 1962 1022
rect 2038 1018 2042 1022
rect 2150 1018 2154 1022
rect 2182 1018 2186 1022
rect 2398 1018 2402 1022
rect 2854 1018 2858 1022
rect 3390 1018 3394 1022
rect 3526 1018 3530 1022
rect 3734 1018 3738 1022
rect 4062 1018 4066 1022
rect 394 1003 398 1007
rect 401 1003 405 1007
rect 1418 1003 1422 1007
rect 1425 1003 1429 1007
rect 2442 1003 2446 1007
rect 2449 1003 2453 1007
rect 3474 1003 3478 1007
rect 3481 1003 3485 1007
rect 30 988 34 992
rect 206 988 210 992
rect 294 988 298 992
rect 438 988 442 992
rect 662 988 666 992
rect 854 988 858 992
rect 886 988 890 992
rect 942 988 946 992
rect 1054 988 1058 992
rect 1094 988 1098 992
rect 1406 988 1410 992
rect 1534 988 1538 992
rect 1574 988 1578 992
rect 1590 988 1594 992
rect 1630 988 1634 992
rect 1806 988 1810 992
rect 1902 988 1906 992
rect 1942 988 1946 992
rect 2126 988 2130 992
rect 2142 988 2146 992
rect 2302 988 2306 992
rect 2582 988 2586 992
rect 2686 988 2690 992
rect 3094 988 3098 992
rect 3542 988 3546 992
rect 3662 988 3666 992
rect 3822 988 3826 992
rect 3998 988 4002 992
rect 4070 988 4074 992
rect 4094 988 4098 992
rect 4142 988 4146 992
rect 4206 988 4210 992
rect 4222 988 4226 992
rect 4270 988 4274 992
rect 4286 988 4290 992
rect 262 978 266 982
rect 614 979 618 983
rect 1990 978 1994 982
rect 3158 978 3162 982
rect 3326 979 3330 983
rect 6 968 10 972
rect 486 968 490 972
rect 1022 968 1026 972
rect 2742 968 2746 972
rect 3846 968 3850 972
rect 4006 968 4010 972
rect 4038 968 4042 972
rect 4062 968 4066 972
rect 4102 968 4106 972
rect 4134 968 4138 972
rect 4198 968 4202 972
rect 4230 968 4234 972
rect 4246 968 4250 972
rect 206 958 210 962
rect 238 958 242 962
rect 254 958 258 962
rect 438 958 442 962
rect 614 956 618 960
rect 694 958 698 962
rect 854 958 858 962
rect 974 958 978 962
rect 982 958 986 962
rect 1174 958 1178 962
rect 1286 958 1290 962
rect 1318 958 1322 962
rect 1326 958 1330 962
rect 1462 958 1466 962
rect 1494 958 1498 962
rect 1718 958 1722 962
rect 1822 958 1826 962
rect 1854 958 1858 962
rect 1886 958 1890 962
rect 2302 958 2306 962
rect 2478 958 2482 962
rect 2622 958 2626 962
rect 2758 958 2762 962
rect 2790 958 2794 962
rect 2862 958 2866 962
rect 3094 958 3098 962
rect 3118 958 3122 962
rect 3166 958 3170 962
rect 3326 956 3330 960
rect 3382 958 3386 962
rect 3494 958 3498 962
rect 3574 958 3578 962
rect 3590 958 3594 962
rect 3606 958 3610 962
rect 3734 958 3738 962
rect 3790 958 3794 962
rect 3990 958 3994 962
rect 4022 958 4026 962
rect 4078 958 4082 962
rect 4086 958 4090 962
rect 4118 958 4122 962
rect 4182 958 4186 962
rect 4214 958 4218 962
rect 4246 958 4250 962
rect 4302 958 4306 962
rect 22 948 26 952
rect 198 948 202 952
rect 238 948 242 952
rect 286 948 290 952
rect 438 948 442 952
rect 526 948 530 952
rect 622 948 626 952
rect 750 948 754 952
rect 902 948 906 952
rect 1030 948 1034 952
rect 1062 948 1066 952
rect 1110 948 1114 952
rect 1134 948 1138 952
rect 1142 948 1146 952
rect 1158 948 1162 952
rect 1190 948 1194 952
rect 1198 948 1202 952
rect 1214 948 1218 952
rect 1222 948 1226 952
rect 1254 948 1258 952
rect 1270 948 1274 952
rect 1302 948 1306 952
rect 1342 948 1346 952
rect 1358 948 1362 952
rect 1366 948 1370 952
rect 1390 948 1394 952
rect 1446 948 1450 952
rect 1478 948 1482 952
rect 1494 948 1498 952
rect 1526 948 1530 952
rect 1558 948 1562 952
rect 1574 948 1578 952
rect 1614 948 1618 952
rect 1670 948 1674 952
rect 1694 948 1698 952
rect 1710 948 1714 952
rect 1758 948 1762 952
rect 1790 948 1794 952
rect 1806 948 1810 952
rect 1846 948 1850 952
rect 1862 948 1866 952
rect 1870 948 1874 952
rect 1902 948 1906 952
rect 1934 948 1938 952
rect 1958 948 1962 952
rect 1974 948 1978 952
rect 1982 948 1986 952
rect 2030 948 2034 952
rect 2054 948 2058 952
rect 2070 948 2074 952
rect 2078 948 2082 952
rect 2102 948 2106 952
rect 2110 948 2114 952
rect 2198 948 2202 952
rect 2326 948 2330 952
rect 2358 948 2362 952
rect 2366 948 2370 952
rect 2406 948 2410 952
rect 2430 948 2434 952
rect 2446 948 2450 952
rect 2478 948 2482 952
rect 2486 948 2490 952
rect 2502 948 2506 952
rect 2518 948 2522 952
rect 2550 948 2554 952
rect 2622 948 2626 952
rect 2670 948 2674 952
rect 2686 948 2690 952
rect 2734 948 2738 952
rect 2774 948 2778 952
rect 2798 948 2802 952
rect 2838 948 2842 952
rect 2878 948 2882 952
rect 2886 948 2890 952
rect 3086 948 3090 952
rect 3134 948 3138 952
rect 3238 948 3242 952
rect 3406 948 3410 952
rect 3422 948 3426 952
rect 3438 948 3442 952
rect 3470 948 3474 952
rect 3502 948 3506 952
rect 3510 948 3514 952
rect 3518 948 3522 952
rect 3590 948 3594 952
rect 3614 948 3618 952
rect 3646 948 3650 952
rect 3702 948 3706 952
rect 3718 948 3722 952
rect 3766 948 3770 952
rect 3798 948 3802 952
rect 3830 948 3834 952
rect 3918 948 3922 952
rect 3934 948 3938 952
rect 3966 948 3970 952
rect 3998 948 4002 952
rect 4030 948 4034 952
rect 4046 948 4050 952
rect 4070 948 4074 952
rect 4094 948 4098 952
rect 4126 948 4130 952
rect 4174 948 4178 952
rect 4190 948 4194 952
rect 4222 948 4226 952
rect 4254 948 4258 952
rect 4286 948 4290 952
rect 4310 948 4314 952
rect 4374 948 4378 952
rect 158 938 162 942
rect 230 938 234 942
rect 390 938 394 942
rect 582 938 586 942
rect 654 938 658 942
rect 670 938 674 942
rect 806 938 810 942
rect 950 938 954 942
rect 998 938 1002 942
rect 1006 938 1010 942
rect 1030 938 1034 942
rect 1062 938 1066 942
rect 1070 938 1074 942
rect 1078 938 1082 942
rect 1150 938 1154 942
rect 1166 938 1170 942
rect 1230 938 1234 942
rect 1262 938 1266 942
rect 1294 938 1298 942
rect 1350 938 1354 942
rect 1438 938 1442 942
rect 1454 938 1458 942
rect 1470 938 1474 942
rect 1542 938 1546 942
rect 1582 938 1586 942
rect 1606 938 1610 942
rect 1638 938 1642 942
rect 1798 938 1802 942
rect 1878 938 1882 942
rect 1910 938 1914 942
rect 2022 938 2026 942
rect 2118 938 2122 942
rect 2134 938 2138 942
rect 2254 938 2258 942
rect 2334 938 2338 942
rect 2350 938 2354 942
rect 2454 938 2458 942
rect 2494 938 2498 942
rect 2526 938 2530 942
rect 2534 938 2538 942
rect 2542 938 2546 942
rect 2590 938 2594 942
rect 2598 938 2602 942
rect 2614 938 2618 942
rect 2662 938 2666 942
rect 2678 938 2682 942
rect 2734 938 2738 942
rect 2742 938 2746 942
rect 2766 938 2770 942
rect 2806 938 2810 942
rect 2822 938 2826 942
rect 2846 938 2850 942
rect 2870 938 2874 942
rect 2902 938 2906 942
rect 2934 938 2938 942
rect 3046 938 3050 942
rect 3126 938 3130 942
rect 3150 938 3154 942
rect 3190 938 3194 942
rect 3197 938 3201 942
rect 3294 938 3298 942
rect 3366 938 3370 942
rect 3398 938 3402 942
rect 3414 938 3418 942
rect 3438 938 3442 942
rect 3446 938 3450 942
rect 3462 938 3466 942
rect 3518 938 3522 942
rect 3550 938 3554 942
rect 3558 938 3562 942
rect 3582 938 3586 942
rect 3622 938 3626 942
rect 3670 938 3674 942
rect 3710 938 3714 942
rect 3742 938 3746 942
rect 3758 938 3762 942
rect 3774 938 3778 942
rect 3806 938 3810 942
rect 3822 938 3826 942
rect 3902 938 3906 942
rect 3910 938 3914 942
rect 3958 938 3962 942
rect 4278 938 4282 942
rect 142 928 146 932
rect 374 928 378 932
rect 566 928 570 932
rect 702 928 706 932
rect 710 928 714 932
rect 790 928 794 932
rect 1094 928 1098 932
rect 1126 928 1130 932
rect 1374 928 1378 932
rect 1430 928 1434 932
rect 1510 928 1514 932
rect 1542 928 1546 932
rect 1598 928 1602 932
rect 1646 928 1650 932
rect 1710 928 1714 932
rect 1718 928 1722 932
rect 1742 928 1746 932
rect 1830 928 1834 932
rect 1918 928 1922 932
rect 1958 928 1962 932
rect 2158 928 2162 932
rect 2238 928 2242 932
rect 2342 928 2346 932
rect 2382 928 2386 932
rect 2390 928 2394 932
rect 2510 928 2514 932
rect 2646 928 2650 932
rect 2710 928 2714 932
rect 2822 928 2826 932
rect 2918 928 2922 932
rect 3030 928 3034 932
rect 3278 928 3282 932
rect 3454 928 3458 932
rect 3638 928 3642 932
rect 3742 928 3746 932
rect 3942 928 3946 932
rect 974 918 978 922
rect 982 918 986 922
rect 1014 918 1018 922
rect 1286 918 1290 922
rect 1318 918 1322 922
rect 1326 918 1330 922
rect 1678 918 1682 922
rect 1774 918 1778 922
rect 1838 918 1842 922
rect 2086 918 2090 922
rect 2374 918 2378 922
rect 2398 918 2402 922
rect 2566 918 2570 922
rect 2606 918 2610 922
rect 2790 918 2794 922
rect 2814 918 2818 922
rect 2950 918 2954 922
rect 3166 918 3170 922
rect 3374 918 3378 922
rect 3390 918 3394 922
rect 3630 918 3634 922
rect 3686 918 3690 922
rect 3750 918 3754 922
rect 3782 918 3786 922
rect 4158 918 4162 922
rect 4326 918 4330 922
rect 4350 918 4354 922
rect 898 903 902 907
rect 905 903 909 907
rect 1930 903 1934 907
rect 1937 903 1941 907
rect 2954 903 2958 907
rect 2961 903 2965 907
rect 3978 903 3982 907
rect 3985 903 3989 907
rect 614 888 618 892
rect 646 888 650 892
rect 790 888 794 892
rect 1006 888 1010 892
rect 1230 888 1234 892
rect 1278 888 1282 892
rect 1334 888 1338 892
rect 1494 888 1498 892
rect 1662 888 1666 892
rect 1758 888 1762 892
rect 2102 888 2106 892
rect 2382 888 2386 892
rect 2446 888 2450 892
rect 2478 888 2482 892
rect 2598 888 2602 892
rect 2662 888 2666 892
rect 2742 888 2746 892
rect 2774 888 2778 892
rect 3054 888 3058 892
rect 3198 888 3202 892
rect 3542 888 3546 892
rect 3726 888 3730 892
rect 3790 888 3794 892
rect 3918 888 3922 892
rect 4054 888 4058 892
rect 4118 888 4122 892
rect 4150 888 4154 892
rect 4182 888 4186 892
rect 4198 888 4202 892
rect 4222 888 4226 892
rect 4254 888 4258 892
rect 4278 888 4282 892
rect 4342 888 4346 892
rect 142 878 146 882
rect 438 878 442 882
rect 694 878 698 882
rect 806 878 810 882
rect 926 878 930 882
rect 1022 878 1026 882
rect 1046 878 1050 882
rect 1134 878 1138 882
rect 1342 878 1346 882
rect 1406 878 1410 882
rect 1430 878 1434 882
rect 1462 878 1466 882
rect 1654 878 1658 882
rect 1702 878 1706 882
rect 1726 878 1730 882
rect 1982 878 1986 882
rect 2070 878 2074 882
rect 2086 878 2090 882
rect 2110 878 2114 882
rect 2118 878 2122 882
rect 2206 878 2210 882
rect 2534 878 2538 882
rect 2590 878 2594 882
rect 2678 878 2682 882
rect 2782 878 2786 882
rect 2870 878 2874 882
rect 2982 878 2986 882
rect 3094 878 3098 882
rect 3110 878 3114 882
rect 3118 878 3122 882
rect 3222 878 3226 882
rect 3310 878 3314 882
rect 3382 878 3386 882
rect 3438 878 3442 882
rect 3622 878 3626 882
rect 3734 878 3738 882
rect 3846 878 3850 882
rect 4158 878 4162 882
rect 4190 878 4194 882
rect 6 868 10 872
rect 30 868 34 872
rect 158 868 162 872
rect 230 868 234 872
rect 262 868 266 872
rect 334 868 338 872
rect 454 868 458 872
rect 558 868 562 872
rect 662 868 666 872
rect 678 868 682 872
rect 742 868 746 872
rect 758 868 762 872
rect 910 868 914 872
rect 1150 868 1154 872
rect 1222 868 1226 872
rect 1262 868 1266 872
rect 1270 868 1274 872
rect 1294 868 1298 872
rect 1326 868 1330 872
rect 1350 868 1354 872
rect 1382 868 1386 872
rect 1454 868 1458 872
rect 1550 868 1554 872
rect 1582 868 1586 872
rect 1590 868 1594 872
rect 1646 868 1650 872
rect 1734 868 1738 872
rect 1782 868 1786 872
rect 1798 868 1802 872
rect 1806 868 1810 872
rect 1822 868 1826 872
rect 1838 868 1842 872
rect 1998 868 2002 872
rect 2222 868 2226 872
rect 2294 868 2298 872
rect 2358 868 2362 872
rect 2366 868 2370 872
rect 2414 868 2418 872
rect 2422 868 2426 872
rect 2470 868 2474 872
rect 2486 868 2490 872
rect 2502 868 2506 872
rect 2518 868 2522 872
rect 2550 868 2554 872
rect 2582 868 2586 872
rect 2606 868 2610 872
rect 2622 868 2626 872
rect 2670 868 2674 872
rect 2694 868 2698 872
rect 2710 868 2714 872
rect 2758 868 2762 872
rect 2766 868 2770 872
rect 2806 868 2810 872
rect 2814 868 2818 872
rect 2822 868 2826 872
rect 2830 868 2834 872
rect 2862 868 2866 872
rect 2894 868 2898 872
rect 2926 868 2930 872
rect 2934 868 2938 872
rect 2966 868 2970 872
rect 3014 868 3018 872
rect 3046 868 3050 872
rect 3078 868 3082 872
rect 3102 868 3106 872
rect 3134 868 3138 872
rect 3190 868 3194 872
rect 3206 868 3210 872
rect 3246 868 3250 872
rect 3254 868 3258 872
rect 3342 868 3346 872
rect 3350 868 3354 872
rect 3398 868 3402 872
rect 3422 868 3426 872
rect 3438 868 3442 872
rect 3454 868 3458 872
rect 3470 868 3474 872
rect 3526 868 3530 872
rect 3638 868 3642 872
rect 3718 868 3722 872
rect 3734 868 3738 872
rect 3766 868 3770 872
rect 3782 868 3786 872
rect 3798 868 3802 872
rect 3814 868 3818 872
rect 3862 868 3866 872
rect 3894 868 3898 872
rect 3902 868 3906 872
rect 4094 868 4098 872
rect 4142 868 4146 872
rect 4158 868 4162 872
rect 4206 868 4210 872
rect 22 858 26 862
rect 46 858 50 862
rect 198 858 202 862
rect 238 858 242 862
rect 454 858 458 862
rect 510 858 514 862
rect 550 858 554 862
rect 630 858 634 862
rect 670 858 674 862
rect 686 858 690 862
rect 718 858 722 862
rect 750 858 754 862
rect 774 858 778 862
rect 798 858 802 862
rect 822 858 826 862
rect 870 858 874 862
rect 1038 858 1042 862
rect 1094 858 1098 862
rect 1206 858 1210 862
rect 1302 858 1306 862
rect 1318 858 1322 862
rect 1350 858 1354 862
rect 1374 858 1378 862
rect 1390 858 1394 862
rect 1454 858 1458 862
rect 1478 858 1482 862
rect 1494 858 1498 862
rect 1510 858 1514 862
rect 1542 858 1546 862
rect 1574 858 1578 862
rect 1638 858 1642 862
rect 1670 858 1674 862
rect 1686 858 1690 862
rect 1710 858 1714 862
rect 1758 858 1762 862
rect 1766 858 1770 862
rect 1790 858 1794 862
rect 1806 858 1810 862
rect 1830 858 1834 862
rect 1846 858 1850 862
rect 1870 858 1874 862
rect 1901 858 1905 862
rect 1942 858 1946 862
rect 2054 858 2058 862
rect 2070 858 2074 862
rect 2094 858 2098 862
rect 2166 858 2170 862
rect 2310 858 2314 862
rect 2406 858 2410 862
rect 2462 858 2466 862
rect 2494 858 2498 862
rect 2510 858 2514 862
rect 2558 858 2562 862
rect 2614 858 2618 862
rect 2630 858 2634 862
rect 2638 858 2642 862
rect 2734 858 2738 862
rect 2798 858 2802 862
rect 2838 858 2842 862
rect 2870 858 2874 862
rect 2918 858 2922 862
rect 2942 858 2946 862
rect 2958 858 2962 862
rect 2990 858 2994 862
rect 3038 858 3042 862
rect 3070 858 3074 862
rect 3142 858 3146 862
rect 3174 858 3178 862
rect 3214 858 3218 862
rect 3238 858 3242 862
rect 3262 858 3266 862
rect 3286 858 3290 862
rect 3334 858 3338 862
rect 3358 858 3362 862
rect 3406 858 3410 862
rect 3414 858 3418 862
rect 3446 858 3450 862
rect 3478 858 3482 862
rect 3502 858 3506 862
rect 3518 858 3522 862
rect 3638 858 3642 862
rect 3678 858 3682 862
rect 3710 858 3714 862
rect 3758 858 3762 862
rect 3774 858 3778 862
rect 3806 858 3810 862
rect 3822 858 3826 862
rect 3838 858 3842 862
rect 3870 858 3874 862
rect 3934 858 3938 862
rect 3974 858 3978 862
rect 4014 858 4018 862
rect 4030 858 4034 862
rect 4046 858 4050 862
rect 4078 858 4082 862
rect 4118 858 4122 862
rect 4134 858 4138 862
rect 4166 858 4170 862
rect 4238 858 4242 862
rect 4270 858 4274 862
rect 4294 858 4298 862
rect 4318 858 4322 862
rect 4358 858 4362 862
rect 62 848 66 852
rect 206 848 210 852
rect 254 848 258 852
rect 486 850 490 854
rect 686 848 690 852
rect 710 848 714 852
rect 766 848 770 852
rect 878 850 882 854
rect 1182 850 1186 854
rect 1246 848 1250 852
rect 1358 848 1362 852
rect 1526 848 1530 852
rect 1558 848 1562 852
rect 1614 848 1618 852
rect 1702 848 1706 852
rect 1774 848 1778 852
rect 2030 850 2034 854
rect 2254 850 2258 854
rect 2302 848 2306 852
rect 2342 848 2346 852
rect 2390 848 2394 852
rect 2438 848 2442 852
rect 2566 848 2570 852
rect 2646 848 2650 852
rect 2654 848 2658 852
rect 2742 848 2746 852
rect 2782 848 2786 852
rect 2870 848 2874 852
rect 2902 848 2906 852
rect 2942 848 2946 852
rect 2990 848 2994 852
rect 3022 848 3026 852
rect 3054 848 3058 852
rect 3222 848 3226 852
rect 3278 848 3282 852
rect 3318 848 3322 852
rect 3334 848 3338 852
rect 3502 848 3506 852
rect 3686 848 3690 852
rect 3742 848 3746 852
rect 3878 848 3882 852
rect 3918 848 3922 852
rect 3926 848 3930 852
rect 3998 848 4002 852
rect 4006 848 4010 852
rect 4062 848 4066 852
rect 4070 848 4074 852
rect 4126 848 4130 852
rect 4302 848 4306 852
rect 4310 848 4314 852
rect 4366 848 4370 852
rect 238 838 242 842
rect 358 838 362 842
rect 726 838 730 842
rect 1238 838 1242 842
rect 1286 838 1290 842
rect 1302 838 1306 842
rect 1598 838 1602 842
rect 2358 838 2362 842
rect 3942 838 3946 842
rect 3966 838 3970 842
rect 4014 838 4018 842
rect 4022 838 4026 842
rect 4046 838 4050 842
rect 4086 838 4090 842
rect 4110 838 4114 842
rect 4286 838 4290 842
rect 4326 838 4330 842
rect 4334 838 4338 842
rect 4350 838 4354 842
rect 486 827 490 831
rect 878 827 882 831
rect 2030 827 2034 831
rect 3086 828 3090 832
rect 3358 828 3362 832
rect 3470 828 3474 832
rect 206 818 210 822
rect 534 818 538 822
rect 718 818 722 822
rect 1038 818 1042 822
rect 1182 818 1186 822
rect 1254 818 1258 822
rect 1574 818 1578 822
rect 1638 818 1642 822
rect 2254 818 2258 822
rect 2326 818 2330 822
rect 2678 818 2682 822
rect 2774 818 2778 822
rect 2838 818 2842 822
rect 3134 818 3138 822
rect 3166 818 3170 822
rect 3310 818 3314 822
rect 3686 818 3690 822
rect 3934 818 3938 822
rect 394 803 398 807
rect 401 803 405 807
rect 1418 803 1422 807
rect 1425 803 1429 807
rect 2442 803 2446 807
rect 2449 803 2453 807
rect 3474 803 3478 807
rect 3481 803 3485 807
rect 30 788 34 792
rect 206 788 210 792
rect 390 788 394 792
rect 574 788 578 792
rect 614 788 618 792
rect 790 788 794 792
rect 934 788 938 792
rect 1022 788 1026 792
rect 1102 788 1106 792
rect 1390 788 1394 792
rect 1406 788 1410 792
rect 1430 788 1434 792
rect 1502 788 1506 792
rect 1534 788 1538 792
rect 1558 788 1562 792
rect 1582 788 1586 792
rect 1670 788 1674 792
rect 1702 788 1706 792
rect 1734 788 1738 792
rect 1806 788 1810 792
rect 1822 788 1826 792
rect 1982 788 1986 792
rect 2046 788 2050 792
rect 2078 788 2082 792
rect 2222 788 2226 792
rect 2366 788 2370 792
rect 2566 788 2570 792
rect 2678 788 2682 792
rect 3054 788 3058 792
rect 3254 788 3258 792
rect 3326 788 3330 792
rect 3470 788 3474 792
rect 3646 788 3650 792
rect 3766 788 3770 792
rect 3862 788 3866 792
rect 3886 788 3890 792
rect 3926 788 3930 792
rect 3958 788 3962 792
rect 4006 788 4010 792
rect 4038 788 4042 792
rect 4062 788 4066 792
rect 4134 788 4138 792
rect 4190 788 4194 792
rect 4230 788 4234 792
rect 4326 788 4330 792
rect 430 778 434 782
rect 1350 779 1354 783
rect 1614 778 1618 782
rect 2806 779 2810 783
rect 3182 779 3186 783
rect 6 768 10 772
rect 310 768 314 772
rect 678 768 682 772
rect 766 768 770 772
rect 1174 768 1178 772
rect 1190 768 1194 772
rect 2598 768 2602 772
rect 2654 768 2658 772
rect 3518 768 3522 772
rect 3822 768 3826 772
rect 3838 768 3842 772
rect 3854 768 3858 772
rect 3878 768 3882 772
rect 3918 768 3922 772
rect 3950 768 3954 772
rect 3998 768 4002 772
rect 4030 768 4034 772
rect 4054 768 4058 772
rect 4126 768 4130 772
rect 4182 768 4186 772
rect 4222 768 4226 772
rect 4278 768 4282 772
rect 4318 768 4322 772
rect 206 758 210 762
rect 326 758 330 762
rect 574 758 578 762
rect 662 758 666 762
rect 726 758 730 762
rect 790 758 794 762
rect 1038 758 1042 762
rect 1158 758 1162 762
rect 1206 758 1210 762
rect 1350 756 1354 760
rect 1518 758 1522 762
rect 1550 758 1554 762
rect 1598 758 1602 762
rect 1686 758 1690 762
rect 1718 758 1722 762
rect 22 748 26 752
rect 198 748 202 752
rect 310 748 314 752
rect 470 748 474 752
rect 598 748 602 752
rect 622 748 626 752
rect 646 748 650 752
rect 670 748 674 752
rect 694 748 698 752
rect 718 748 722 752
rect 726 748 730 752
rect 742 748 746 752
rect 894 748 898 752
rect 1086 748 1090 752
rect 1118 748 1122 752
rect 1150 748 1154 752
rect 1174 748 1178 752
rect 1198 748 1202 752
rect 1262 748 1266 752
rect 1374 748 1378 752
rect 1454 748 1458 752
rect 1470 748 1474 752
rect 1486 748 1490 752
rect 1502 748 1506 752
rect 1518 748 1522 752
rect 1582 748 1586 752
rect 1622 748 1626 752
rect 1662 748 1666 752
rect 1670 748 1674 752
rect 1702 748 1706 752
rect 1734 748 1738 752
rect 1766 758 1770 762
rect 1790 758 1794 762
rect 1950 758 1954 762
rect 2014 758 2018 762
rect 2030 758 2034 762
rect 2062 758 2066 762
rect 2222 758 2226 762
rect 2438 758 2442 762
rect 2494 758 2498 762
rect 2574 758 2578 762
rect 2582 758 2586 762
rect 2598 758 2602 762
rect 2638 758 2642 762
rect 2806 756 2810 760
rect 2886 758 2890 762
rect 2902 758 2906 762
rect 2942 758 2946 762
rect 2958 758 2962 762
rect 2982 758 2986 762
rect 3182 756 3186 760
rect 3470 758 3474 762
rect 3590 758 3594 762
rect 3598 758 3602 762
rect 3694 758 3698 762
rect 3742 758 3746 762
rect 3798 758 3802 762
rect 3806 758 3810 762
rect 3838 758 3842 762
rect 3910 758 3914 762
rect 3934 758 3938 762
rect 3966 758 3970 762
rect 4014 758 4018 762
rect 4070 758 4074 762
rect 4110 758 4114 762
rect 4198 758 4202 762
rect 4206 758 4210 762
rect 4302 758 4306 762
rect 1782 748 1786 752
rect 1806 748 1810 752
rect 1822 748 1826 752
rect 1846 748 1850 752
rect 1886 748 1890 752
rect 1934 748 1938 752
rect 1966 748 1970 752
rect 1982 748 1986 752
rect 2014 748 2018 752
rect 2046 748 2050 752
rect 2222 748 2226 752
rect 2246 748 2250 752
rect 2302 748 2306 752
rect 2350 748 2354 752
rect 2406 748 2410 752
rect 2422 748 2426 752
rect 2446 748 2450 752
rect 2462 748 2466 752
rect 2478 748 2482 752
rect 2510 748 2514 752
rect 2526 748 2530 752
rect 2630 748 2634 752
rect 2654 748 2658 752
rect 2814 748 2818 752
rect 2846 748 2850 752
rect 2878 748 2882 752
rect 2902 748 2906 752
rect 2918 748 2922 752
rect 2998 748 3002 752
rect 3038 748 3042 752
rect 3094 748 3098 752
rect 3222 748 3226 752
rect 3278 748 3282 752
rect 3294 748 3298 752
rect 3462 748 3466 752
rect 3518 748 3522 752
rect 3566 748 3570 752
rect 3614 748 3618 752
rect 3630 748 3634 752
rect 3662 748 3666 752
rect 3726 748 3730 752
rect 3750 748 3754 752
rect 3814 748 3818 752
rect 3846 748 3850 752
rect 3886 748 3890 752
rect 3910 748 3914 752
rect 3942 748 3946 752
rect 3990 748 3994 752
rect 4022 748 4026 752
rect 4062 748 4066 752
rect 4102 748 4106 752
rect 4118 748 4122 752
rect 4166 748 4170 752
rect 4190 748 4194 752
rect 4214 748 4218 752
rect 4238 748 4242 752
rect 4294 748 4298 752
rect 4310 748 4314 752
rect 4358 748 4362 752
rect 4390 748 4394 752
rect 158 738 162 742
rect 230 738 234 742
rect 294 738 298 742
rect 302 738 306 742
rect 334 738 338 742
rect 526 738 530 742
rect 654 738 658 742
rect 718 738 722 742
rect 838 738 842 742
rect 966 738 970 742
rect 1078 738 1082 742
rect 1142 738 1146 742
rect 1158 738 1162 742
rect 1221 738 1225 742
rect 1318 738 1322 742
rect 1462 738 1466 742
rect 1478 738 1482 742
rect 1494 738 1498 742
rect 1526 738 1530 742
rect 1574 738 1578 742
rect 1630 738 1634 742
rect 1646 738 1650 742
rect 1662 738 1666 742
rect 1694 738 1698 742
rect 1726 738 1730 742
rect 1814 738 1818 742
rect 1894 738 1898 742
rect 1926 738 1930 742
rect 1974 738 1978 742
rect 2006 738 2010 742
rect 2038 738 2042 742
rect 2174 738 2178 742
rect 2270 738 2274 742
rect 2294 738 2298 742
rect 2358 738 2362 742
rect 2382 738 2386 742
rect 2398 738 2402 742
rect 2414 738 2418 742
rect 2470 738 2474 742
rect 2502 738 2506 742
rect 2518 738 2522 742
rect 2534 738 2538 742
rect 2558 738 2562 742
rect 2598 738 2602 742
rect 2622 738 2626 742
rect 2670 738 2674 742
rect 2774 738 2778 742
rect 2854 738 2858 742
rect 2878 738 2882 742
rect 2910 738 2914 742
rect 2918 738 2922 742
rect 2934 738 2938 742
rect 2966 738 2970 742
rect 3006 738 3010 742
rect 3046 738 3050 742
rect 3150 738 3154 742
rect 3246 738 3250 742
rect 3270 738 3274 742
rect 3286 738 3290 742
rect 3302 738 3306 742
rect 3422 738 3426 742
rect 3510 738 3514 742
rect 3558 738 3562 742
rect 3574 738 3578 742
rect 3622 738 3626 742
rect 3710 738 3714 742
rect 3718 738 3722 742
rect 3782 738 3786 742
rect 3798 738 3802 742
rect 4254 738 4258 742
rect 142 728 146 732
rect 510 728 514 732
rect 766 728 770 732
rect 854 728 858 732
rect 1062 728 1066 732
rect 1126 728 1130 732
rect 1302 728 1306 732
rect 1398 728 1402 732
rect 1430 728 1434 732
rect 1446 728 1450 732
rect 1566 728 1570 732
rect 1606 728 1610 732
rect 1838 728 1842 732
rect 1870 728 1874 732
rect 1910 728 1914 732
rect 1998 728 2002 732
rect 2158 728 2162 732
rect 2278 728 2282 732
rect 2486 728 2490 732
rect 2550 728 2554 732
rect 2606 728 2610 732
rect 2758 728 2762 732
rect 3014 728 3018 732
rect 3134 728 3138 732
rect 3222 728 3226 732
rect 3238 728 3242 732
rect 3406 728 3410 732
rect 3542 728 3546 732
rect 3582 728 3586 732
rect 3742 728 3746 732
rect 1038 718 1042 722
rect 1102 718 1106 722
rect 1134 718 1138 722
rect 1166 718 1170 722
rect 1638 718 1642 722
rect 1854 718 1858 722
rect 1878 718 1882 722
rect 1902 718 1906 722
rect 1918 718 1922 722
rect 2286 718 2290 722
rect 2318 718 2322 722
rect 2334 718 2338 722
rect 2398 718 2402 722
rect 2542 718 2546 722
rect 2862 718 2866 722
rect 2974 718 2978 722
rect 2982 718 2986 722
rect 3022 718 3026 722
rect 3310 718 3314 722
rect 3598 718 3602 722
rect 3678 718 3682 722
rect 3702 718 3706 722
rect 3766 718 3770 722
rect 4086 718 4090 722
rect 4150 718 4154 722
rect 4342 718 4346 722
rect 4374 718 4378 722
rect 898 703 902 707
rect 905 703 909 707
rect 1930 703 1934 707
rect 1937 703 1941 707
rect 2954 703 2958 707
rect 2961 703 2965 707
rect 3978 703 3982 707
rect 3985 703 3989 707
rect 214 688 218 692
rect 734 688 738 692
rect 766 688 770 692
rect 878 688 882 692
rect 926 688 930 692
rect 958 688 962 692
rect 1238 688 1242 692
rect 1510 688 1514 692
rect 1526 688 1530 692
rect 1622 688 1626 692
rect 1686 688 1690 692
rect 1846 688 1850 692
rect 1998 688 2002 692
rect 2366 688 2370 692
rect 2582 688 2586 692
rect 2590 688 2594 692
rect 2622 688 2626 692
rect 2646 688 2650 692
rect 2870 688 2874 692
rect 2926 688 2930 692
rect 3206 688 3210 692
rect 3742 688 3746 692
rect 3910 688 3914 692
rect 3998 688 4002 692
rect 4158 688 4162 692
rect 4214 688 4218 692
rect 4246 688 4250 692
rect 118 678 122 682
rect 366 678 370 682
rect 630 678 634 682
rect 782 678 786 682
rect 1126 678 1130 682
rect 1558 678 1562 682
rect 1654 678 1658 682
rect 1766 678 1770 682
rect 1774 678 1778 682
rect 1910 678 1914 682
rect 1974 678 1978 682
rect 2078 678 2082 682
rect 2182 678 2186 682
rect 2230 678 2234 682
rect 2294 678 2298 682
rect 2358 678 2362 682
rect 2390 678 2394 682
rect 2486 678 2490 682
rect 2630 678 2634 682
rect 2846 678 2850 682
rect 2878 678 2882 682
rect 3030 678 3034 682
rect 3110 678 3114 682
rect 3198 678 3202 682
rect 3246 678 3250 682
rect 3270 678 3274 682
rect 3302 678 3306 682
rect 3334 678 3338 682
rect 3342 678 3346 682
rect 3358 678 3362 682
rect 3590 678 3594 682
rect 3686 678 3690 682
rect 3774 678 3778 682
rect 3782 678 3786 682
rect 3854 678 3858 682
rect 3886 678 3890 682
rect 4126 678 4130 682
rect 4166 678 4170 682
rect 4238 678 4242 682
rect 4390 678 4394 682
rect 134 668 138 672
rect 270 668 274 672
rect 382 668 386 672
rect 470 668 474 672
rect 534 668 538 672
rect 646 668 650 672
rect 822 668 826 672
rect 982 668 986 672
rect 998 668 1002 672
rect 1110 668 1114 672
rect 1230 668 1234 672
rect 1246 668 1250 672
rect 1270 668 1274 672
rect 1286 668 1290 672
rect 1350 668 1354 672
rect 1358 668 1362 672
rect 1374 668 1378 672
rect 1454 668 1458 672
rect 1470 668 1474 672
rect 1486 668 1490 672
rect 1518 668 1522 672
rect 1550 668 1554 672
rect 1614 668 1618 672
rect 1646 668 1650 672
rect 1678 668 1682 672
rect 1710 668 1714 672
rect 1718 668 1722 672
rect 1734 668 1738 672
rect 1750 668 1754 672
rect 2094 668 2098 672
rect 2190 668 2194 672
rect 2222 668 2226 672
rect 2254 668 2258 672
rect 2286 668 2290 672
rect 2310 668 2314 672
rect 2502 668 2506 672
rect 2574 668 2578 672
rect 2614 668 2618 672
rect 2654 668 2658 672
rect 2662 668 2666 672
rect 2718 668 2722 672
rect 2734 668 2738 672
rect 2750 668 2754 672
rect 2766 668 2770 672
rect 2790 668 2794 672
rect 2830 668 2834 672
rect 2854 668 2858 672
rect 2918 668 2922 672
rect 2966 668 2970 672
rect 3014 668 3018 672
rect 3126 668 3130 672
rect 3214 668 3218 672
rect 3294 668 3298 672
rect 3326 668 3330 672
rect 3414 668 3418 672
rect 3422 668 3426 672
rect 3510 668 3514 672
rect 3542 668 3546 672
rect 3550 668 3554 672
rect 3566 668 3570 672
rect 3630 668 3634 672
rect 3678 668 3682 672
rect 3694 668 3698 672
rect 3718 668 3722 672
rect 3750 668 3754 672
rect 3798 668 3802 672
rect 3830 668 3834 672
rect 3846 668 3850 672
rect 3870 668 3874 672
rect 4150 668 4154 672
rect 4166 668 4170 672
rect 4254 668 4258 672
rect 4278 668 4282 672
rect 4350 668 4354 672
rect 4358 668 4362 672
rect 182 658 186 662
rect 326 658 330 662
rect 438 658 442 662
rect 590 658 594 662
rect 702 658 706 662
rect 718 658 722 662
rect 750 658 754 662
rect 806 658 810 662
rect 838 658 842 662
rect 862 658 866 662
rect 886 658 890 662
rect 934 658 938 662
rect 974 658 978 662
rect 1006 658 1010 662
rect 1030 658 1034 662
rect 1110 658 1114 662
rect 1214 658 1218 662
rect 1254 658 1258 662
rect 1262 658 1266 662
rect 1294 658 1298 662
rect 1318 658 1322 662
rect 1350 658 1354 662
rect 1390 658 1394 662
rect 1422 658 1426 662
rect 1430 658 1434 662
rect 1438 658 1442 662
rect 1462 658 1466 662
rect 1494 658 1498 662
rect 1526 658 1530 662
rect 1606 658 1610 662
rect 1622 658 1626 662
rect 1670 658 1674 662
rect 1686 658 1690 662
rect 1702 658 1706 662
rect 1726 658 1730 662
rect 1750 658 1754 662
rect 1790 658 1794 662
rect 1822 658 1826 662
rect 1838 658 1842 662
rect 1862 658 1866 662
rect 1870 658 1874 662
rect 1902 658 1906 662
rect 1942 658 1946 662
rect 2094 658 2098 662
rect 2166 658 2170 662
rect 2198 658 2202 662
rect 2214 658 2218 662
rect 2278 658 2282 662
rect 2286 658 2290 662
rect 2318 658 2322 662
rect 2326 658 2330 662
rect 2390 658 2394 662
rect 2502 658 2506 662
rect 2614 658 2618 662
rect 2670 658 2674 662
rect 2710 658 2714 662
rect 2726 658 2730 662
rect 2758 658 2762 662
rect 2798 658 2802 662
rect 2822 658 2826 662
rect 2838 658 2842 662
rect 2854 658 2858 662
rect 2886 658 2890 662
rect 2910 658 2914 662
rect 2942 658 2946 662
rect 2950 658 2954 662
rect 2958 658 2962 662
rect 3006 658 3010 662
rect 3070 658 3074 662
rect 3222 658 3226 662
rect 3230 658 3234 662
rect 3254 658 3258 662
rect 3358 658 3362 662
rect 3382 658 3386 662
rect 3406 658 3410 662
rect 3478 658 3482 662
rect 3502 658 3506 662
rect 3534 658 3538 662
rect 3574 658 3578 662
rect 3606 658 3610 662
rect 3670 658 3674 662
rect 3726 658 3730 662
rect 3758 658 3762 662
rect 3806 658 3810 662
rect 3846 658 3850 662
rect 3878 658 3882 662
rect 3910 658 3914 662
rect 3942 658 3946 662
rect 3998 658 4002 662
rect 4022 658 4026 662
rect 4038 658 4042 662
rect 4062 658 4066 662
rect 4086 658 4090 662
rect 4102 658 4106 662
rect 4126 658 4130 662
rect 4142 658 4146 662
rect 4198 658 4202 662
rect 4214 658 4218 662
rect 4262 658 4266 662
rect 4278 658 4282 662
rect 4310 658 4314 662
rect 4334 658 4338 662
rect 4366 658 4370 662
rect 182 648 186 652
rect 414 650 418 654
rect 694 648 698 652
rect 822 648 826 652
rect 830 648 834 652
rect 998 648 1002 652
rect 1038 648 1042 652
rect 1078 650 1082 654
rect 1286 648 1290 652
rect 1334 648 1338 652
rect 1382 648 1386 652
rect 1478 648 1482 652
rect 1510 648 1514 652
rect 1590 648 1594 652
rect 1742 648 1746 652
rect 2142 648 2146 652
rect 2174 648 2178 652
rect 2230 648 2234 652
rect 2334 648 2338 652
rect 2350 648 2354 652
rect 2534 650 2538 654
rect 2590 648 2594 652
rect 2638 648 2642 652
rect 2686 648 2690 652
rect 2694 648 2698 652
rect 2782 648 2786 652
rect 2798 648 2802 652
rect 2814 648 2818 652
rect 2990 648 2994 652
rect 3006 648 3010 652
rect 3174 648 3178 652
rect 3390 648 3394 652
rect 3406 648 3410 652
rect 3494 648 3498 652
rect 3534 648 3538 652
rect 3614 648 3618 652
rect 3646 648 3650 652
rect 3654 648 3658 652
rect 3742 648 3746 652
rect 3774 648 3778 652
rect 3822 648 3826 652
rect 3830 648 3834 652
rect 3902 648 3906 652
rect 3934 648 3938 652
rect 4006 648 4010 652
rect 4014 648 4018 652
rect 4070 648 4074 652
rect 4078 648 4082 652
rect 4134 648 4138 652
rect 4206 648 4210 652
rect 4270 648 4274 652
rect 4302 648 4306 652
rect 6 638 10 642
rect 846 638 850 642
rect 1022 638 1026 642
rect 1310 638 1314 642
rect 2206 638 2210 642
rect 2262 638 2266 642
rect 3630 638 3634 642
rect 3918 638 3922 642
rect 3950 638 3954 642
rect 3974 638 3978 642
rect 3990 638 3994 642
rect 3998 638 4002 642
rect 4022 638 4026 642
rect 4030 638 4034 642
rect 4054 638 4058 642
rect 4062 638 4066 642
rect 4094 638 4098 642
rect 4118 638 4122 642
rect 4214 638 4218 642
rect 4286 638 4290 642
rect 4318 638 4322 642
rect 1014 628 1018 632
rect 1078 627 1082 631
rect 3806 628 3810 632
rect 4310 628 4314 632
rect 182 618 186 622
rect 214 618 218 622
rect 286 618 290 622
rect 414 618 418 622
rect 550 618 554 622
rect 694 618 698 622
rect 790 618 794 622
rect 838 618 842 622
rect 1206 618 1210 622
rect 1302 618 1306 622
rect 1406 618 1410 622
rect 1782 618 1786 622
rect 1806 618 1810 622
rect 1886 618 1890 622
rect 1934 618 1938 622
rect 1958 618 1962 622
rect 1982 618 1986 622
rect 2142 618 2146 622
rect 2534 618 2538 622
rect 2622 618 2626 622
rect 2670 618 2674 622
rect 2710 618 2714 622
rect 2750 618 2754 622
rect 3174 618 3178 622
rect 3230 618 3234 622
rect 3254 618 3258 622
rect 3278 618 3282 622
rect 3310 618 3314 622
rect 3350 618 3354 622
rect 3374 618 3378 622
rect 3430 618 3434 622
rect 3566 618 3570 622
rect 3710 618 3714 622
rect 3790 618 3794 622
rect 3894 618 3898 622
rect 4390 618 4394 622
rect 394 603 398 607
rect 401 603 405 607
rect 1418 603 1422 607
rect 1425 603 1429 607
rect 2442 603 2446 607
rect 2449 603 2453 607
rect 3474 603 3478 607
rect 3481 603 3485 607
rect 166 588 170 592
rect 198 588 202 592
rect 558 588 562 592
rect 614 588 618 592
rect 758 588 762 592
rect 854 588 858 592
rect 934 588 938 592
rect 1078 588 1082 592
rect 1310 588 1314 592
rect 1350 588 1354 592
rect 1462 588 1466 592
rect 1486 588 1490 592
rect 1518 588 1522 592
rect 1582 588 1586 592
rect 1646 588 1650 592
rect 1726 588 1730 592
rect 1766 588 1770 592
rect 1814 588 1818 592
rect 1878 588 1882 592
rect 2166 588 2170 592
rect 2438 588 2442 592
rect 2582 588 2586 592
rect 2894 588 2898 592
rect 3342 588 3346 592
rect 3486 588 3490 592
rect 3638 588 3642 592
rect 3710 588 3714 592
rect 3926 588 3930 592
rect 3966 588 3970 592
rect 4006 588 4010 592
rect 4022 588 4026 592
rect 4070 588 4074 592
rect 4118 588 4122 592
rect 4182 588 4186 592
rect 4214 588 4218 592
rect 4254 588 4258 592
rect 4278 588 4282 592
rect 4358 588 4362 592
rect 4374 588 4378 592
rect 246 579 250 583
rect 1182 579 1186 583
rect 3022 579 3026 583
rect 3070 578 3074 582
rect 4102 578 4106 582
rect 1382 568 1386 572
rect 1790 568 1794 572
rect 1918 568 1922 572
rect 3126 568 3130 572
rect 3918 568 3922 572
rect 3950 568 3954 572
rect 3966 568 3970 572
rect 4030 568 4034 572
rect 4062 568 4066 572
rect 4094 568 4098 572
rect 4126 568 4130 572
rect 4158 568 4162 572
rect 4190 568 4194 572
rect 4222 568 4226 572
rect 4246 568 4250 572
rect 4286 568 4290 572
rect 4318 568 4322 572
rect 4382 568 4386 572
rect 246 556 250 560
rect 406 558 410 562
rect 758 558 762 562
rect 806 558 810 562
rect 814 558 818 562
rect 934 558 938 562
rect 1094 558 1098 562
rect 1158 558 1162 562
rect 78 548 82 552
rect 150 548 154 552
rect 174 548 178 552
rect 182 548 186 552
rect 230 548 234 552
rect 422 548 426 552
rect 438 548 442 552
rect 542 548 546 552
rect 582 548 586 552
rect 710 548 714 552
rect 742 548 746 552
rect 790 548 794 552
rect 838 548 842 552
rect 870 548 874 552
rect 1038 548 1042 552
rect 1142 548 1146 552
rect 1182 556 1186 560
rect 1414 558 1418 562
rect 1446 558 1450 562
rect 1502 558 1506 562
rect 1534 558 1538 562
rect 1630 558 1634 562
rect 1662 558 1666 562
rect 1694 558 1698 562
rect 1990 558 1994 562
rect 2038 558 2042 562
rect 2182 558 2186 562
rect 2222 558 2226 562
rect 2238 558 2242 562
rect 1270 548 1274 552
rect 1326 548 1330 552
rect 1334 548 1338 552
rect 1358 548 1362 552
rect 1382 548 1386 552
rect 1430 548 1434 552
rect 1454 548 1458 552
rect 1486 548 1490 552
rect 1510 548 1514 552
rect 1542 548 1546 552
rect 1558 548 1562 552
rect 1574 548 1578 552
rect 1590 548 1594 552
rect 1614 548 1618 552
rect 1622 548 1626 552
rect 1638 548 1642 552
rect 1678 548 1682 552
rect 1710 548 1714 552
rect 1726 548 1730 552
rect 1742 548 1746 552
rect 1766 548 1770 552
rect 1806 548 1810 552
rect 1846 548 1850 552
rect 1878 548 1882 552
rect 1902 548 1906 552
rect 1934 548 1938 552
rect 1942 548 1946 552
rect 1974 548 1978 552
rect 1998 548 2002 552
rect 2086 548 2090 552
rect 2118 548 2122 552
rect 2150 548 2154 552
rect 2158 548 2162 552
rect 2206 548 2210 552
rect 2222 548 2226 552
rect 2254 548 2258 552
rect 2278 558 2282 562
rect 2390 558 2394 562
rect 2406 558 2410 562
rect 2582 558 2586 562
rect 2606 558 2610 562
rect 2702 558 2706 562
rect 2710 558 2714 562
rect 2814 558 2818 562
rect 3022 556 3026 560
rect 3206 558 3210 562
rect 3326 558 3330 562
rect 3486 558 3490 562
rect 3590 558 3594 562
rect 3726 558 3730 562
rect 3782 558 3786 562
rect 3806 558 3810 562
rect 3830 558 3834 562
rect 3870 558 3874 562
rect 3894 558 3898 562
rect 3902 558 3906 562
rect 3934 558 3938 562
rect 3982 558 3986 562
rect 4014 558 4018 562
rect 4046 558 4050 562
rect 4078 558 4082 562
rect 4110 558 4114 562
rect 4142 558 4146 562
rect 4174 558 4178 562
rect 4206 558 4210 562
rect 4262 558 4266 562
rect 4270 558 4274 562
rect 4302 558 4306 562
rect 4334 558 4338 562
rect 4366 558 4370 562
rect 2294 548 2298 552
rect 2326 548 2330 552
rect 2358 548 2362 552
rect 2390 548 2394 552
rect 2478 548 2482 552
rect 2582 548 2586 552
rect 2646 548 2650 552
rect 2734 548 2738 552
rect 2782 548 2786 552
rect 2822 548 2826 552
rect 2934 548 2938 552
rect 3038 548 3042 552
rect 3110 548 3114 552
rect 3126 548 3130 552
rect 3174 548 3178 552
rect 3190 548 3194 552
rect 3214 548 3218 552
rect 3246 548 3250 552
rect 3310 548 3314 552
rect 3470 548 3474 552
rect 3534 548 3538 552
rect 3582 548 3586 552
rect 3654 548 3658 552
rect 3750 548 3754 552
rect 3910 548 3914 552
rect 3942 548 3946 552
rect 3990 548 3994 552
rect 4022 548 4026 552
rect 4054 548 4058 552
rect 4086 548 4090 552
rect 4118 548 4122 552
rect 4126 548 4130 552
rect 4150 548 4154 552
rect 4166 548 4170 552
rect 4182 548 4186 552
rect 4214 548 4218 552
rect 4254 548 4258 552
rect 4278 548 4282 552
rect 4310 548 4314 552
rect 4342 548 4346 552
rect 4374 548 4378 552
rect 6 538 10 542
rect 142 538 146 542
rect 278 538 282 542
rect 430 538 434 542
rect 470 538 474 542
rect 534 538 538 542
rect 574 538 578 542
rect 710 538 714 542
rect 782 538 786 542
rect 798 538 802 542
rect 830 538 834 542
rect 982 538 986 542
rect 1118 538 1122 542
rect 1214 538 1218 542
rect 1374 538 1378 542
rect 1422 538 1426 542
rect 1438 538 1442 542
rect 1478 538 1482 542
rect 1510 538 1514 542
rect 1566 538 1570 542
rect 1598 538 1602 542
rect 1606 538 1610 542
rect 1638 538 1642 542
rect 1670 538 1674 542
rect 1966 538 1970 542
rect 1982 538 1986 542
rect 2022 538 2026 542
rect 2046 538 2050 542
rect 2158 538 2162 542
rect 2214 538 2218 542
rect 2246 538 2250 542
rect 2262 538 2266 542
rect 2350 538 2354 542
rect 2382 538 2386 542
rect 2534 538 2538 542
rect 2622 538 2626 542
rect 2670 540 2674 544
rect 2678 538 2682 542
rect 2686 538 2690 542
rect 2726 538 2730 542
rect 2790 538 2794 542
rect 2798 538 2802 542
rect 2854 538 2858 542
rect 2990 538 2994 542
rect 3062 538 3066 542
rect 3086 538 3090 542
rect 3094 538 3098 542
rect 3110 538 3114 542
rect 3118 538 3122 542
rect 3166 538 3170 542
rect 3182 538 3186 542
rect 3222 538 3226 542
rect 3254 538 3258 542
rect 3270 538 3274 542
rect 3310 538 3314 542
rect 3438 538 3442 542
rect 3518 538 3522 542
rect 3574 538 3578 542
rect 3614 538 3618 542
rect 3646 538 3650 542
rect 3686 538 3690 542
rect 3742 538 3746 542
rect 3798 538 3802 542
rect 3822 538 3826 542
rect 3846 538 3850 542
rect 3878 538 3882 542
rect 294 528 298 532
rect 694 528 698 532
rect 998 528 1002 532
rect 1086 528 1090 532
rect 1230 528 1234 532
rect 1470 528 1474 532
rect 1558 528 1562 532
rect 1758 528 1762 532
rect 1782 528 1786 532
rect 1790 528 1794 532
rect 1822 528 1826 532
rect 1830 528 1834 532
rect 1846 528 1850 532
rect 1870 528 1874 532
rect 1878 528 1882 532
rect 1894 528 1898 532
rect 2014 528 2018 532
rect 2054 528 2058 532
rect 2134 528 2138 532
rect 2190 528 2194 532
rect 2206 528 2210 532
rect 2302 528 2306 532
rect 2342 528 2346 532
rect 2518 528 2522 532
rect 2630 528 2634 532
rect 2750 528 2754 532
rect 2846 528 2850 532
rect 2974 528 2978 532
rect 3150 528 3154 532
rect 3230 528 3234 532
rect 3238 528 3242 532
rect 3422 528 3426 532
rect 3558 528 3562 532
rect 62 518 66 522
rect 406 518 410 522
rect 454 518 458 522
rect 598 518 602 522
rect 814 518 818 522
rect 886 518 890 522
rect 1126 518 1130 522
rect 1310 518 1314 522
rect 2006 518 2010 522
rect 2030 518 2034 522
rect 2102 518 2106 522
rect 2334 518 2338 522
rect 2374 518 2378 522
rect 2606 518 2610 522
rect 2638 518 2642 522
rect 2654 518 2658 522
rect 2694 518 2698 522
rect 2710 518 2714 522
rect 2766 518 2770 522
rect 2814 518 2818 522
rect 2838 518 2842 522
rect 2878 518 2882 522
rect 3070 518 3074 522
rect 3206 518 3210 522
rect 3262 518 3266 522
rect 3318 518 3322 522
rect 3550 518 3554 522
rect 3598 518 3602 522
rect 3670 518 3674 522
rect 3734 518 3738 522
rect 3766 518 3770 522
rect 3790 518 3794 522
rect 3814 518 3818 522
rect 3830 518 3834 522
rect 3862 518 3866 522
rect 3894 518 3898 522
rect 898 503 902 507
rect 905 503 909 507
rect 1930 503 1934 507
rect 1937 503 1941 507
rect 2954 503 2958 507
rect 2961 503 2965 507
rect 3978 503 3982 507
rect 3985 503 3989 507
rect 758 488 762 492
rect 1110 488 1114 492
rect 1462 488 1466 492
rect 1494 488 1498 492
rect 1518 488 1522 492
rect 1558 488 1562 492
rect 1574 488 1578 492
rect 1598 488 1602 492
rect 1622 488 1626 492
rect 1654 488 1658 492
rect 1710 488 1714 492
rect 1758 488 1762 492
rect 1910 488 1914 492
rect 2422 488 2426 492
rect 2790 488 2794 492
rect 2854 488 2858 492
rect 3110 488 3114 492
rect 3302 488 3306 492
rect 3550 488 3554 492
rect 3998 488 4002 492
rect 4190 488 4194 492
rect 4246 488 4250 492
rect 4286 488 4290 492
rect 4374 488 4378 492
rect 118 478 122 482
rect 286 478 290 482
rect 654 478 658 482
rect 862 478 866 482
rect 974 478 978 482
rect 1046 478 1050 482
rect 1054 478 1058 482
rect 1270 478 1274 482
rect 1486 478 1490 482
rect 1526 478 1530 482
rect 1566 478 1570 482
rect 1606 478 1610 482
rect 1630 478 1634 482
rect 1750 478 1754 482
rect 1990 478 1994 482
rect 2254 478 2258 482
rect 2550 478 2554 482
rect 2558 478 2562 482
rect 2686 478 2690 482
rect 2934 478 2938 482
rect 3102 478 3106 482
rect 3158 478 3162 482
rect 3406 478 3410 482
rect 3534 478 3538 482
rect 3614 478 3618 482
rect 3846 478 3850 482
rect 3878 478 3882 482
rect 3918 478 3922 482
rect 4198 478 4202 482
rect 4294 478 4298 482
rect 4310 478 4314 482
rect 134 468 138 472
rect 270 468 274 472
rect 398 468 402 472
rect 470 468 474 472
rect 670 468 674 472
rect 878 468 882 472
rect 982 468 986 472
rect 1102 468 1106 472
rect 1126 468 1130 472
rect 1134 468 1138 472
rect 1166 468 1170 472
rect 1254 468 1258 472
rect 1398 468 1402 472
rect 1414 468 1418 472
rect 1454 468 1458 472
rect 1470 468 1474 472
rect 1534 468 1538 472
rect 1638 468 1642 472
rect 1686 468 1690 472
rect 1742 468 1746 472
rect 1766 468 1770 472
rect 1814 466 1818 470
rect 1822 468 1826 472
rect 1830 468 1834 472
rect 1878 468 1882 472
rect 2006 468 2010 472
rect 2078 468 2082 472
rect 2094 468 2098 472
rect 2134 468 2138 472
rect 2142 468 2146 472
rect 2270 468 2274 472
rect 2366 468 2370 472
rect 2374 468 2378 472
rect 2390 468 2394 472
rect 2478 468 2482 472
rect 2486 468 2490 472
rect 2518 468 2522 472
rect 2542 468 2546 472
rect 2702 468 2706 472
rect 2774 468 2778 472
rect 2798 468 2802 472
rect 2806 468 2810 472
rect 2950 468 2954 472
rect 3046 468 3050 472
rect 3062 468 3066 472
rect 3094 468 3098 472
rect 3118 468 3122 472
rect 3142 468 3146 472
rect 3174 468 3178 472
rect 3182 468 3186 472
rect 3190 468 3194 472
rect 3206 468 3210 472
rect 3238 468 3242 472
rect 3310 468 3314 472
rect 3422 468 3426 472
rect 3518 468 3522 472
rect 3566 468 3570 472
rect 3582 468 3586 472
rect 3630 468 3634 472
rect 3646 468 3650 472
rect 3702 468 3706 472
rect 3710 468 3714 472
rect 3750 468 3754 472
rect 3758 468 3762 472
rect 3790 468 3794 472
rect 3822 468 3826 472
rect 3862 468 3866 472
rect 3886 468 3890 472
rect 3934 468 3938 472
rect 4006 468 4010 472
rect 4062 468 4066 472
rect 4158 468 4162 472
rect 4182 468 4186 472
rect 4222 468 4226 472
rect 4278 468 4282 472
rect 182 458 186 462
rect 230 458 234 462
rect 326 458 330 462
rect 542 458 546 462
rect 718 458 722 462
rect 742 458 746 462
rect 822 458 826 462
rect 990 458 994 462
rect 1022 458 1026 462
rect 1078 458 1082 462
rect 1094 458 1098 462
rect 1134 458 1138 462
rect 1142 458 1146 462
rect 1214 458 1218 462
rect 1390 458 1394 462
rect 1406 458 1410 462
rect 1446 458 1450 462
rect 1486 458 1490 462
rect 1510 458 1514 462
rect 1542 458 1546 462
rect 1582 458 1586 462
rect 1590 458 1594 462
rect 1614 458 1618 462
rect 1670 458 1674 462
rect 1694 458 1698 462
rect 1750 458 1754 462
rect 1774 458 1778 462
rect 1790 458 1794 462
rect 1838 458 1842 462
rect 1870 458 1874 462
rect 2038 458 2042 462
rect 2134 458 2138 462
rect 2318 458 2322 462
rect 2358 458 2362 462
rect 2366 458 2370 462
rect 2406 458 2410 462
rect 2454 458 2458 462
rect 2478 458 2482 462
rect 2510 458 2514 462
rect 2526 458 2530 462
rect 2534 458 2538 462
rect 2590 458 2594 462
rect 2646 458 2650 462
rect 2742 458 2746 462
rect 2774 458 2778 462
rect 2814 458 2818 462
rect 2822 458 2826 462
rect 2894 458 2898 462
rect 3054 458 3058 462
rect 3070 458 3074 462
rect 3094 458 3098 462
rect 3134 458 3138 462
rect 3166 458 3170 462
rect 3198 458 3202 462
rect 3230 458 3234 462
rect 3246 458 3250 462
rect 3270 458 3274 462
rect 3286 458 3290 462
rect 3422 458 3426 462
rect 3510 458 3514 462
rect 3542 458 3546 462
rect 3574 458 3578 462
rect 3590 458 3594 462
rect 3638 458 3642 462
rect 3646 458 3650 462
rect 3694 458 3698 462
rect 3726 458 3730 462
rect 3782 458 3786 462
rect 3798 458 3802 462
rect 3822 458 3826 462
rect 3838 458 3842 462
rect 3854 458 3858 462
rect 3870 458 3874 462
rect 3894 458 3898 462
rect 3902 458 3906 462
rect 3942 458 3946 462
rect 3958 458 3962 462
rect 4022 458 4026 462
rect 4038 458 4042 462
rect 4062 458 4066 462
rect 4086 458 4090 462
rect 4102 458 4106 462
rect 4126 458 4130 462
rect 4158 458 4162 462
rect 4174 458 4178 462
rect 4214 458 4218 462
rect 4246 458 4250 462
rect 4270 458 4274 462
rect 166 450 170 454
rect 222 448 226 452
rect 702 450 706 454
rect 910 450 914 454
rect 990 448 994 452
rect 1014 448 1018 452
rect 1086 448 1090 452
rect 1182 448 1186 452
rect 1222 450 1226 454
rect 1438 448 1442 452
rect 1558 448 1562 452
rect 1654 448 1658 452
rect 1710 448 1714 452
rect 1718 448 1722 452
rect 1734 448 1738 452
rect 1790 448 1794 452
rect 1854 448 1858 452
rect 2054 448 2058 452
rect 2110 448 2114 452
rect 2158 448 2162 452
rect 2302 450 2306 454
rect 2342 448 2346 452
rect 2358 448 2362 452
rect 2398 448 2402 452
rect 2510 448 2514 452
rect 2574 448 2578 452
rect 2750 448 2754 452
rect 2822 448 2826 452
rect 2838 448 2842 452
rect 2982 450 2986 454
rect 3038 448 3042 452
rect 3070 448 3074 452
rect 3158 448 3162 452
rect 3262 448 3266 452
rect 3270 448 3274 452
rect 3470 448 3474 452
rect 3590 448 3594 452
rect 3678 448 3682 452
rect 3814 448 3818 452
rect 3950 448 3954 452
rect 3982 448 3986 452
rect 4014 448 4018 452
rect 4070 448 4074 452
rect 4078 448 4082 452
rect 4134 448 4138 452
rect 4166 448 4170 452
rect 4206 448 4210 452
rect 4262 448 4266 452
rect 4302 448 4306 452
rect 4342 458 4346 462
rect 4374 458 4378 462
rect 4334 448 4338 452
rect 4366 448 4370 452
rect 6 438 10 442
rect 558 438 562 442
rect 1030 438 1034 442
rect 1070 438 1074 442
rect 1142 438 1146 442
rect 2126 438 2130 442
rect 2142 438 2146 442
rect 2166 438 2170 442
rect 2606 438 2610 442
rect 3966 438 3970 442
rect 4030 438 4034 442
rect 4054 438 4058 442
rect 4094 438 4098 442
rect 4118 438 4122 442
rect 4150 438 4154 442
rect 4222 438 4226 442
rect 4246 438 4250 442
rect 4310 438 4314 442
rect 4318 438 4322 442
rect 4334 438 4338 442
rect 4382 438 4386 442
rect 366 428 370 432
rect 910 427 914 431
rect 1222 427 1226 431
rect 1646 428 1650 432
rect 2302 427 2306 431
rect 2982 427 2986 431
rect 4126 428 4130 432
rect 4342 428 4346 432
rect 166 418 170 422
rect 222 418 226 422
rect 526 418 530 422
rect 574 418 578 422
rect 702 418 706 422
rect 782 418 786 422
rect 966 418 970 422
rect 1062 418 1066 422
rect 1350 418 1354 422
rect 1374 418 1378 422
rect 1774 418 1778 422
rect 2054 418 2058 422
rect 2086 418 2090 422
rect 2102 418 2106 422
rect 2750 418 2754 422
rect 3214 418 3218 422
rect 3246 418 3250 422
rect 3470 418 3474 422
rect 3654 418 3658 422
rect 3718 418 3722 422
rect 3798 418 3802 422
rect 3982 418 3986 422
rect 394 403 398 407
rect 401 403 405 407
rect 1418 403 1422 407
rect 1425 403 1429 407
rect 2442 403 2446 407
rect 2449 403 2453 407
rect 3474 403 3478 407
rect 3481 403 3485 407
rect 86 388 90 392
rect 254 388 258 392
rect 486 388 490 392
rect 862 388 866 392
rect 1126 388 1130 392
rect 1406 388 1410 392
rect 1646 388 1650 392
rect 1670 388 1674 392
rect 1814 388 1818 392
rect 2030 388 2034 392
rect 2174 388 2178 392
rect 2238 388 2242 392
rect 2766 388 2770 392
rect 2910 388 2914 392
rect 3094 388 3098 392
rect 3438 388 3442 392
rect 4006 388 4010 392
rect 4150 388 4154 392
rect 4182 388 4186 392
rect 4214 388 4218 392
rect 4246 388 4250 392
rect 4278 388 4282 392
rect 4310 388 4314 392
rect 4358 388 4362 392
rect 358 379 362 383
rect 894 368 898 372
rect 1190 378 1194 382
rect 1566 378 1570 382
rect 3222 379 3226 383
rect 3566 379 3570 383
rect 950 368 954 372
rect 1070 368 1074 372
rect 1198 368 1202 372
rect 1310 368 1314 372
rect 1502 368 1506 372
rect 2518 368 2522 372
rect 2574 368 2578 372
rect 3806 368 3810 372
rect 3854 368 3858 372
rect 4190 368 4194 372
rect 4222 368 4226 372
rect 4254 368 4258 372
rect 4286 368 4290 372
rect 4318 368 4322 372
rect 4350 368 4354 372
rect 254 358 258 362
rect 358 356 362 360
rect 558 358 562 362
rect 614 358 618 362
rect 862 358 866 362
rect 926 358 930 362
rect 974 358 978 362
rect 1014 358 1018 362
rect 1038 358 1042 362
rect 1054 358 1058 362
rect 1142 358 1146 362
rect 1182 358 1186 362
rect 1238 358 1242 362
rect 1254 358 1258 362
rect 1286 358 1290 362
rect 1350 358 1354 362
rect 1478 358 1482 362
rect 1518 358 1522 362
rect 1814 358 1818 362
rect 1846 358 1850 362
rect 1950 358 1954 362
rect 2174 358 2178 362
rect 2286 358 2290 362
rect 2318 358 2322 362
rect 2350 358 2354 362
rect 2502 358 2506 362
rect 2534 358 2538 362
rect 2582 358 2586 362
rect 2638 358 2642 362
rect 2702 358 2706 362
rect 2758 358 2762 362
rect 2910 358 2914 362
rect 2982 358 2986 362
rect 2998 358 3002 362
rect 3078 358 3082 362
rect 3222 356 3226 360
rect 3278 358 3282 362
rect 3294 358 3298 362
rect 3334 358 3338 362
rect 3566 356 3570 360
rect 3630 358 3634 362
rect 3670 358 3674 362
rect 3838 358 3842 362
rect 3870 358 3874 362
rect 4150 358 4154 362
rect 4174 358 4178 362
rect 4206 358 4210 362
rect 4238 358 4242 362
rect 4270 358 4274 362
rect 4302 358 4306 362
rect 4334 358 4338 362
rect 30 348 34 352
rect 109 348 113 352
rect 150 348 154 352
rect 254 348 258 352
rect 302 348 306 352
rect 342 348 346 352
rect 518 348 522 352
rect 582 348 586 352
rect 622 348 626 352
rect 646 348 650 352
rect 678 348 682 352
rect 758 348 762 352
rect 846 348 850 352
rect 894 348 898 352
rect 942 348 946 352
rect 974 348 978 352
rect 1022 348 1026 352
rect 1062 348 1066 352
rect 1118 348 1122 352
rect 1126 348 1130 352
rect 1142 348 1146 352
rect 1190 348 1194 352
rect 1230 348 1234 352
rect 1238 348 1242 352
rect 1262 348 1266 352
rect 1294 348 1298 352
rect 1318 348 1322 352
rect 1350 348 1354 352
rect 1398 348 1402 352
rect 1422 348 1426 352
rect 1430 348 1434 352
rect 1454 348 1458 352
rect 1486 348 1490 352
rect 1510 348 1514 352
rect 1526 348 1530 352
rect 1590 348 1594 352
rect 1798 348 1802 352
rect 1838 348 1842 352
rect 1870 348 1874 352
rect 2006 348 2010 352
rect 2070 348 2074 352
rect 2206 348 2210 352
rect 2254 348 2258 352
rect 2270 348 2274 352
rect 2286 348 2290 352
rect 2334 348 2338 352
rect 2366 348 2370 352
rect 2414 348 2418 352
rect 2430 348 2434 352
rect 2470 348 2474 352
rect 2486 348 2490 352
rect 2550 348 2554 352
rect 2606 348 2610 352
rect 2630 348 2634 352
rect 2654 348 2658 352
rect 2694 348 2698 352
rect 2718 348 2722 352
rect 2734 348 2738 352
rect 2806 348 2810 352
rect 2894 348 2898 352
rect 2902 348 2906 352
rect 2998 348 3002 352
rect 3014 348 3018 352
rect 3046 348 3050 352
rect 3062 348 3066 352
rect 3238 348 3242 352
rect 3294 348 3298 352
rect 3302 348 3306 352
rect 3334 348 3338 352
rect 3342 348 3346 352
rect 3374 348 3378 352
rect 3382 348 3386 352
rect 3478 348 3482 352
rect 3614 348 3618 352
rect 3638 348 3642 352
rect 3662 348 3666 352
rect 3710 348 3714 352
rect 3774 348 3778 352
rect 3830 348 3834 352
rect 3854 348 3858 352
rect 3886 348 3890 352
rect 3902 348 3906 352
rect 3934 348 3938 352
rect 3942 348 3946 352
rect 3982 348 3986 352
rect 4134 348 4138 352
rect 4182 348 4186 352
rect 4214 348 4218 352
rect 4246 348 4250 352
rect 4278 348 4282 352
rect 4310 348 4314 352
rect 4342 348 4346 352
rect 6 338 10 342
rect 30 338 34 342
rect 206 338 210 342
rect 278 338 282 342
rect 390 338 394 342
rect 526 338 530 342
rect 590 338 594 342
rect 814 338 818 342
rect 886 338 890 342
rect 966 338 970 342
rect 998 338 1002 342
rect 1110 338 1114 342
rect 1270 338 1274 342
rect 1286 338 1290 342
rect 1334 338 1338 342
rect 1382 338 1386 342
rect 1462 338 1466 342
rect 1478 338 1482 342
rect 1558 338 1562 342
rect 1590 338 1594 342
rect 1766 338 1770 342
rect 1846 338 1850 342
rect 1862 338 1866 342
rect 1942 338 1946 342
rect 1982 338 1986 342
rect 2014 338 2018 342
rect 2126 338 2130 342
rect 2198 338 2202 342
rect 2246 338 2250 342
rect 2262 338 2266 342
rect 2278 338 2282 342
rect 2310 338 2314 342
rect 2342 338 2346 342
rect 2358 338 2362 342
rect 2374 338 2378 342
rect 2398 338 2402 342
rect 2454 338 2458 342
rect 2462 338 2466 342
rect 2494 338 2498 342
rect 2526 338 2530 342
rect 2558 338 2562 342
rect 2566 338 2570 342
rect 2598 338 2602 342
rect 2622 338 2626 342
rect 2662 338 2666 342
rect 2686 338 2690 342
rect 2734 338 2738 342
rect 2862 338 2866 342
rect 2966 338 2970 342
rect 2974 338 2978 342
rect 3006 338 3010 342
rect 3022 338 3026 342
rect 3038 338 3042 342
rect 3054 338 3058 342
rect 3086 338 3090 342
rect 3190 338 3194 342
rect 3262 338 3266 342
rect 3270 338 3274 342
rect 3302 338 3306 342
rect 3310 338 3314 342
rect 3350 338 3354 342
rect 3366 338 3370 342
rect 3422 338 3426 342
rect 3534 338 3538 342
rect 3606 338 3610 342
rect 3670 338 3674 342
rect 3718 338 3722 342
rect 3750 338 3754 342
rect 3822 338 3826 342
rect 3862 338 3866 342
rect 3894 338 3898 342
rect 3910 338 3914 342
rect 3926 338 3930 342
rect 3950 338 3954 342
rect 3966 338 3970 342
rect 4102 338 4106 342
rect 190 328 194 332
rect 406 328 410 332
rect 694 328 698 332
rect 798 328 802 332
rect 1086 328 1090 332
rect 1222 328 1226 332
rect 1302 328 1306 332
rect 1750 328 1754 332
rect 1886 328 1890 332
rect 2110 328 2114 332
rect 2230 328 2234 332
rect 2382 328 2386 332
rect 2606 328 2610 332
rect 2638 328 2642 332
rect 2670 328 2674 332
rect 2702 328 2706 332
rect 2846 328 2850 332
rect 2942 328 2946 332
rect 3174 328 3178 332
rect 3518 328 3522 332
rect 3734 328 3738 332
rect 3766 328 3770 332
rect 3806 328 3810 332
rect 4086 328 4090 332
rect 502 318 506 322
rect 534 318 538 322
rect 614 318 618 322
rect 638 318 642 322
rect 662 318 666 322
rect 718 318 722 322
rect 1166 318 1170 322
rect 1494 318 1498 322
rect 1646 318 1650 322
rect 1990 318 1994 322
rect 2222 318 2226 322
rect 2238 318 2242 322
rect 2390 318 2394 322
rect 2486 318 2490 322
rect 2582 318 2586 322
rect 2678 318 2682 322
rect 2750 318 2754 322
rect 2934 318 2938 322
rect 3030 318 3034 322
rect 3358 318 3362 322
rect 3398 318 3402 322
rect 3646 318 3650 322
rect 3758 318 3762 322
rect 3790 318 3794 322
rect 3870 318 3874 322
rect 3918 318 3922 322
rect 3958 318 3962 322
rect 898 303 902 307
rect 905 303 909 307
rect 1930 303 1934 307
rect 1937 303 1941 307
rect 2954 303 2958 307
rect 2961 303 2965 307
rect 3978 303 3982 307
rect 3985 303 3989 307
rect 766 288 770 292
rect 1254 288 1258 292
rect 1542 288 1546 292
rect 1606 288 1610 292
rect 1814 288 1818 292
rect 2294 288 2298 292
rect 2326 288 2330 292
rect 2606 288 2610 292
rect 2814 288 2818 292
rect 3158 288 3162 292
rect 3334 288 3338 292
rect 3382 288 3386 292
rect 3502 288 3506 292
rect 3606 288 3610 292
rect 3630 288 3634 292
rect 3798 288 3802 292
rect 4046 288 4050 292
rect 4278 288 4282 292
rect 4350 288 4354 292
rect 94 278 98 282
rect 262 278 266 282
rect 518 278 522 282
rect 686 278 690 282
rect 838 278 842 282
rect 1046 278 1050 282
rect 1150 278 1154 282
rect 1510 278 1514 282
rect 1710 278 1714 282
rect 1926 278 1930 282
rect 2086 278 2090 282
rect 2094 278 2098 282
rect 2366 278 2370 282
rect 2566 278 2570 282
rect 2686 278 2690 282
rect 2942 278 2946 282
rect 3238 278 3242 282
rect 3414 278 3418 282
rect 3526 278 3530 282
rect 3614 278 3618 282
rect 3982 278 3986 282
rect 4198 278 4202 282
rect 110 268 114 272
rect 246 268 250 272
rect 382 268 386 272
rect 534 268 538 272
rect 670 268 674 272
rect 806 268 810 272
rect 822 268 826 272
rect 854 268 858 272
rect 926 268 930 272
rect 1030 268 1034 272
rect 1134 268 1138 272
rect 1174 268 1178 272
rect 1206 268 1210 272
rect 1230 268 1234 272
rect 1238 268 1242 272
rect 1270 268 1274 272
rect 1286 268 1290 272
rect 1334 268 1338 272
rect 1366 268 1370 272
rect 1382 268 1386 272
rect 1446 268 1450 272
rect 1470 268 1474 272
rect 1486 268 1490 272
rect 1494 268 1498 272
rect 1526 268 1530 272
rect 1550 268 1554 272
rect 1566 268 1570 272
rect 1582 268 1586 272
rect 1614 268 1618 272
rect 1622 268 1626 272
rect 1726 268 1730 272
rect 1806 268 1810 272
rect 1822 268 1826 272
rect 1942 268 1946 272
rect 2030 268 2034 272
rect 2062 268 2066 272
rect 2102 268 2106 272
rect 2126 268 2130 272
rect 2158 268 2162 272
rect 2166 268 2170 272
rect 2198 268 2202 272
rect 2246 268 2250 272
rect 2254 268 2258 272
rect 2302 268 2306 272
rect 2310 268 2314 272
rect 2374 268 2378 272
rect 2446 268 2450 272
rect 2486 268 2490 272
rect 2494 268 2498 272
rect 2526 268 2530 272
rect 2534 268 2538 272
rect 2590 268 2594 272
rect 2702 268 2706 272
rect 2798 268 2802 272
rect 2806 268 2810 272
rect 2846 268 2850 272
rect 2958 268 2962 272
rect 3070 268 3074 272
rect 3078 268 3082 272
rect 3118 268 3122 272
rect 3134 268 3138 272
rect 3254 268 3258 272
rect 3326 268 3330 272
rect 3494 268 3498 272
rect 3542 268 3546 272
rect 3558 268 3562 272
rect 3574 268 3578 272
rect 3598 268 3602 272
rect 3622 268 3626 272
rect 3662 268 3666 272
rect 3678 268 3682 272
rect 3726 268 3730 272
rect 3758 268 3762 272
rect 3766 268 3770 272
rect 3790 268 3794 272
rect 150 258 154 262
rect 166 258 170 262
rect 198 258 202 262
rect 374 258 378 262
rect 406 258 410 262
rect 534 258 538 262
rect 582 258 586 262
rect 630 258 634 262
rect 782 258 786 262
rect 814 258 818 262
rect 830 258 834 262
rect 862 258 866 262
rect 894 258 898 262
rect 942 258 946 262
rect 958 258 962 262
rect 982 258 986 262
rect 1086 258 1090 262
rect 1166 258 1170 262
rect 1214 258 1218 262
rect 1262 258 1266 262
rect 1294 258 1298 262
rect 1310 258 1314 262
rect 1358 258 1362 262
rect 1390 258 1394 262
rect 1414 258 1418 262
rect 3814 266 3818 270
rect 3854 268 3858 272
rect 3870 268 3874 272
rect 3886 268 3890 272
rect 3926 268 3930 272
rect 3934 268 3938 272
rect 3950 268 3954 272
rect 3998 268 4002 272
rect 4014 268 4018 272
rect 4070 268 4074 272
rect 4086 268 4090 272
rect 4102 268 4106 272
rect 4182 268 4186 272
rect 4286 268 4290 272
rect 1494 258 1498 262
rect 1534 258 1538 262
rect 1558 258 1562 262
rect 1598 258 1602 262
rect 1670 258 1674 262
rect 1782 258 1786 262
rect 1798 258 1802 262
rect 1830 258 1834 262
rect 1886 258 1890 262
rect 1998 258 2002 262
rect 2038 258 2042 262
rect 2118 258 2122 262
rect 2150 258 2154 262
rect 2158 258 2162 262
rect 2254 258 2258 262
rect 2278 258 2282 262
rect 2350 258 2354 262
rect 2382 258 2386 262
rect 2430 258 2434 262
rect 2462 258 2466 262
rect 2478 258 2482 262
rect 2502 258 2506 262
rect 2518 258 2522 262
rect 2542 258 2546 262
rect 2590 258 2594 262
rect 2646 258 2650 262
rect 2742 258 2746 262
rect 2782 258 2786 262
rect 2790 258 2794 262
rect 2830 258 2834 262
rect 2838 258 2842 262
rect 2902 258 2906 262
rect 2958 258 2962 262
rect 3046 258 3050 262
rect 3062 258 3066 262
rect 3086 258 3090 262
rect 3094 258 3098 262
rect 3110 258 3114 262
rect 3126 258 3130 262
rect 3142 258 3146 262
rect 3302 258 3306 262
rect 3350 258 3354 262
rect 3366 258 3370 262
rect 3406 258 3410 262
rect 3438 258 3442 262
rect 3486 258 3490 262
rect 3518 258 3522 262
rect 3550 258 3554 262
rect 3566 258 3570 262
rect 3590 258 3594 262
rect 3662 258 3666 262
rect 3702 258 3706 262
rect 3718 258 3722 262
rect 3750 258 3754 262
rect 3774 258 3778 262
rect 3846 258 3850 262
rect 3862 258 3866 262
rect 3894 258 3898 262
rect 3902 258 3906 262
rect 3918 258 3922 262
rect 3942 258 3946 262
rect 4006 258 4010 262
rect 4022 258 4026 262
rect 4038 258 4042 262
rect 4062 258 4066 262
rect 4078 258 4082 262
rect 4110 258 4114 262
rect 4126 258 4130 262
rect 4134 258 4138 262
rect 158 248 162 252
rect 214 250 218 254
rect 358 248 362 252
rect 566 250 570 254
rect 638 250 642 254
rect 830 248 834 252
rect 878 248 882 252
rect 886 248 890 252
rect 958 248 962 252
rect 998 250 1002 254
rect 1182 248 1186 252
rect 1198 248 1202 252
rect 1206 248 1210 252
rect 1286 248 1290 252
rect 1350 248 1354 252
rect 1382 248 1386 252
rect 1422 248 1426 252
rect 1462 248 1466 252
rect 1470 248 1474 252
rect 1534 248 1538 252
rect 1598 248 1602 252
rect 1774 248 1778 252
rect 1974 250 1978 254
rect 2086 248 2090 252
rect 2102 248 2106 252
rect 2134 248 2138 252
rect 2222 248 2226 252
rect 2286 248 2290 252
rect 2334 248 2338 252
rect 2414 248 2418 252
rect 2430 248 2434 252
rect 2462 248 2466 252
rect 2518 248 2522 252
rect 2750 248 2754 252
rect 2774 248 2778 252
rect 2822 248 2826 252
rect 2862 248 2866 252
rect 2990 250 2994 254
rect 3046 248 3050 252
rect 3102 248 3106 252
rect 3286 250 3290 254
rect 3366 248 3370 252
rect 3582 248 3586 252
rect 3638 248 3642 252
rect 3702 248 3706 252
rect 3718 248 3722 252
rect 3734 248 3738 252
rect 3790 248 3794 252
rect 3830 248 3834 252
rect 3902 248 3906 252
rect 3958 248 3962 252
rect 4038 248 4042 252
rect 4046 248 4050 252
rect 4150 250 4154 254
rect 862 238 866 242
rect 894 238 898 242
rect 902 238 906 242
rect 1190 238 1194 242
rect 1254 238 1258 242
rect 1318 238 1322 242
rect 1446 238 1450 242
rect 2150 238 2154 242
rect 3974 238 3978 242
rect 566 227 570 231
rect 638 227 642 231
rect 998 227 1002 231
rect 2038 228 2042 232
rect 3286 227 3290 231
rect 4150 227 4154 231
rect 14 218 18 222
rect 158 218 162 222
rect 214 218 218 222
rect 342 218 346 222
rect 374 218 378 222
rect 422 218 426 222
rect 438 218 442 222
rect 798 218 802 222
rect 1126 218 1130 222
rect 1302 218 1306 222
rect 1398 218 1402 222
rect 1478 218 1482 222
rect 1582 218 1586 222
rect 1774 218 1778 222
rect 1846 218 1850 222
rect 1974 218 1978 222
rect 2174 218 2178 222
rect 2398 218 2402 222
rect 2542 218 2546 222
rect 2750 218 2754 222
rect 2814 218 2818 222
rect 2990 218 2994 222
rect 3454 218 3458 222
rect 3654 218 3658 222
rect 3750 218 3754 222
rect 3870 218 3874 222
rect 4086 218 4090 222
rect 394 203 398 207
rect 401 203 405 207
rect 1418 203 1422 207
rect 1425 203 1429 207
rect 2442 203 2446 207
rect 2449 203 2453 207
rect 3474 203 3478 207
rect 3481 203 3485 207
rect 62 188 66 192
rect 310 188 314 192
rect 870 188 874 192
rect 894 188 898 192
rect 1118 188 1122 192
rect 1246 188 1250 192
rect 1790 188 1794 192
rect 1854 188 1858 192
rect 2222 188 2226 192
rect 2238 188 2242 192
rect 2262 188 2266 192
rect 2806 188 2810 192
rect 2950 188 2954 192
rect 2990 188 2994 192
rect 3110 188 3114 192
rect 3134 188 3138 192
rect 3206 188 3210 192
rect 3350 188 3354 192
rect 3606 188 3610 192
rect 3638 188 3642 192
rect 3998 188 4002 192
rect 4030 188 4034 192
rect 4174 188 4178 192
rect 4286 188 4290 192
rect 4334 188 4338 192
rect 4366 188 4370 192
rect 182 179 186 183
rect 526 179 530 183
rect 726 179 730 183
rect 1086 178 1090 182
rect 830 168 834 172
rect 902 168 906 172
rect 950 168 954 172
rect 958 168 962 172
rect 1006 168 1010 172
rect 1094 168 1098 172
rect 1326 178 1330 182
rect 1582 178 1586 182
rect 2014 178 2018 182
rect 2390 179 2394 183
rect 2614 178 2618 182
rect 3766 179 3770 183
rect 1158 168 1162 172
rect 1230 168 1234 172
rect 1262 168 1266 172
rect 1398 168 1402 172
rect 1494 168 1498 172
rect 2126 168 2130 172
rect 3462 168 3466 172
rect 4206 168 4210 172
rect 182 156 186 160
rect 526 156 530 160
rect 726 156 730 160
rect 790 158 794 162
rect 846 158 850 162
rect 886 158 890 162
rect 934 158 938 162
rect 974 158 978 162
rect 990 158 994 162
rect 1022 158 1026 162
rect 1038 158 1042 162
rect 1054 158 1058 162
rect 1078 158 1082 162
rect 1142 158 1146 162
rect 1214 158 1218 162
rect 1222 158 1226 162
rect 1278 158 1282 162
rect 1310 158 1314 162
rect 1342 158 1346 162
rect 1414 158 1418 162
rect 1462 158 1466 162
rect 1510 158 1514 162
rect 1534 158 1538 162
rect 1790 158 1794 162
rect 1958 158 1962 162
rect 2078 158 2082 162
rect 2086 158 2090 162
rect 2142 158 2146 162
rect 166 148 170 152
rect 342 148 346 152
rect 534 148 538 152
rect 638 148 642 152
rect 806 148 810 152
rect 830 148 834 152
rect 854 148 858 152
rect 894 148 898 152
rect 942 148 946 152
rect 974 148 978 152
rect 1006 148 1010 152
rect 1038 148 1042 152
rect 1086 148 1090 152
rect 1118 148 1122 152
rect 1150 148 1154 152
rect 1198 148 1202 152
rect 1238 148 1242 152
rect 1262 148 1266 152
rect 1286 148 1290 152
rect 1318 148 1322 152
rect 1350 148 1354 152
rect 1382 148 1386 152
rect 1406 148 1410 152
rect 1438 148 1442 152
rect 1470 148 1474 152
rect 1494 148 1498 152
rect 1534 148 1538 152
rect 1558 148 1562 152
rect 1590 148 1594 152
rect 1598 148 1602 152
rect 1614 148 1618 152
rect 1630 148 1634 152
rect 1782 148 1786 152
rect 1830 148 1834 152
rect 1910 148 1914 152
rect 1926 148 1930 152
rect 1974 148 1978 152
rect 2022 148 2026 152
rect 2038 148 2042 152
rect 2054 148 2058 152
rect 2070 148 2074 152
rect 2086 148 2090 152
rect 2102 148 2106 152
rect 2126 148 2130 152
rect 2174 158 2178 162
rect 2390 156 2394 160
rect 2534 158 2538 162
rect 2702 158 2706 162
rect 2750 158 2754 162
rect 2190 148 2194 152
rect 2206 148 2210 152
rect 2230 148 2234 152
rect 2398 148 2402 152
rect 2462 148 2466 152
rect 2494 148 2498 152
rect 2534 148 2538 152
rect 2550 148 2554 152
rect 2566 148 2570 152
rect 2614 148 2618 152
rect 2630 148 2634 152
rect 2662 148 2666 152
rect 2694 148 2698 152
rect 2718 148 2722 152
rect 2806 158 2810 162
rect 3350 158 3354 162
rect 3374 158 3378 162
rect 3606 158 3610 162
rect 3614 158 3618 162
rect 2774 148 2778 152
rect 2910 148 2914 152
rect 3054 148 3058 152
rect 3246 148 3250 152
rect 3334 148 3338 152
rect 3390 148 3394 152
rect 3406 148 3410 152
rect 3502 148 3506 152
rect 3766 156 3770 160
rect 3830 158 3834 162
rect 3902 158 3906 162
rect 3918 158 3922 162
rect 4174 158 4178 162
rect 4270 158 4274 162
rect 4358 158 4362 162
rect 3734 148 3738 152
rect 3774 148 3778 152
rect 3814 148 3818 152
rect 3838 148 3842 152
rect 3854 148 3858 152
rect 3878 148 3882 152
rect 3894 148 3898 152
rect 3918 148 3922 152
rect 3934 148 3938 152
rect 3966 148 3970 152
rect 4014 148 4018 152
rect 4070 148 4074 152
rect 4126 148 4130 152
rect 4286 148 4290 152
rect 4318 148 4322 152
rect 4350 148 4354 152
rect 6 138 10 142
rect 78 138 82 142
rect 142 138 146 142
rect 214 138 218 142
rect 494 138 498 142
rect 694 138 698 142
rect 814 138 818 142
rect 822 138 826 142
rect 966 138 970 142
rect 998 138 1002 142
rect 1030 138 1034 142
rect 1070 138 1074 142
rect 1110 138 1114 142
rect 1190 138 1194 142
rect 1254 138 1258 142
rect 1286 138 1290 142
rect 1302 138 1306 142
rect 1318 138 1322 142
rect 1358 138 1362 142
rect 1374 138 1378 142
rect 1382 138 1386 142
rect 1446 138 1450 142
rect 1462 138 1466 142
rect 1526 138 1530 142
rect 1550 138 1554 142
rect 1566 138 1570 142
rect 1582 138 1586 142
rect 1606 138 1610 142
rect 1622 138 1626 142
rect 1645 138 1649 142
rect 1742 138 1746 142
rect 1814 138 1818 142
rect 1862 138 1866 142
rect 1902 138 1906 142
rect 1918 138 1922 142
rect 1950 138 1954 142
rect 1966 138 1970 142
rect 2030 138 2034 142
rect 2054 138 2058 142
rect 2110 138 2114 142
rect 2118 138 2122 142
rect 2150 138 2154 142
rect 2198 138 2202 142
rect 2358 138 2362 142
rect 2430 138 2434 142
rect 2454 138 2458 142
rect 2470 138 2474 142
rect 2558 138 2562 142
rect 2574 138 2578 142
rect 2622 138 2626 142
rect 2638 138 2642 142
rect 2654 138 2658 142
rect 2726 138 2730 142
rect 2734 138 2738 142
rect 2766 138 2770 142
rect 2782 138 2786 142
rect 2854 138 2858 142
rect 3190 138 3194 142
rect 3302 138 3306 142
rect 3398 138 3402 142
rect 3414 138 3418 142
rect 3430 138 3434 142
rect 3558 138 3562 142
rect 3734 138 3738 142
rect 3806 138 3810 142
rect 3846 138 3850 142
rect 3886 138 3890 142
rect 3926 138 3930 142
rect 3942 138 3946 142
rect 3950 138 3954 142
rect 3958 138 3962 142
rect 3966 138 3970 142
rect 4126 138 4130 142
rect 4262 138 4266 142
rect 4302 138 4306 142
rect 4374 138 4378 142
rect 230 128 234 132
rect 478 128 482 132
rect 678 128 682 132
rect 854 128 858 132
rect 870 128 874 132
rect 878 128 882 132
rect 1062 128 1066 132
rect 1174 128 1178 132
rect 1374 128 1378 132
rect 1726 128 1730 132
rect 1998 128 2002 132
rect 2006 128 2010 132
rect 2046 128 2050 132
rect 2342 128 2346 132
rect 2478 128 2482 132
rect 2502 128 2506 132
rect 2590 128 2594 132
rect 2678 128 2682 132
rect 2870 128 2874 132
rect 3286 128 3290 132
rect 3430 128 3434 132
rect 3542 128 3546 132
rect 3718 128 3722 132
rect 3862 128 3866 132
rect 4110 128 4114 132
rect 4302 128 4306 132
rect 326 118 330 122
rect 350 118 354 122
rect 566 118 570 122
rect 766 118 770 122
rect 1214 118 1218 122
rect 1478 118 1482 122
rect 2158 118 2162 122
rect 2638 118 2642 122
rect 3374 118 3378 122
rect 3830 118 3834 122
rect 4310 118 4314 122
rect 4054 108 4058 112
rect 898 103 902 107
rect 905 103 909 107
rect 1930 103 1934 107
rect 1937 103 1941 107
rect 2954 103 2958 107
rect 2961 103 2965 107
rect 3978 103 3982 107
rect 3985 103 3989 107
rect 310 88 314 92
rect 830 88 834 92
rect 1134 88 1138 92
rect 1334 88 1338 92
rect 1390 88 1394 92
rect 1406 88 1410 92
rect 1598 88 1602 92
rect 1622 88 1626 92
rect 1798 88 1802 92
rect 2046 88 2050 92
rect 2118 88 2122 92
rect 2142 88 2146 92
rect 2174 88 2178 92
rect 2254 88 2258 92
rect 2286 88 2290 92
rect 2318 88 2322 92
rect 2350 88 2354 92
rect 2382 88 2386 92
rect 2406 88 2410 92
rect 2790 88 2794 92
rect 3278 88 3282 92
rect 3350 88 3354 92
rect 3702 88 3706 92
rect 3902 88 3906 92
rect 4038 88 4042 92
rect 4086 88 4090 92
rect 4174 88 4178 92
rect 4214 88 4218 92
rect 4262 88 4266 92
rect 4294 88 4298 92
rect 4334 88 4338 92
rect 4358 88 4362 92
rect 142 78 146 82
rect 526 78 530 82
rect 750 78 754 82
rect 1110 78 1114 82
rect 1142 78 1146 82
rect 1230 78 1234 82
rect 1518 78 1522 82
rect 1702 78 1706 82
rect 1878 78 1882 82
rect 2014 78 2018 82
rect 2190 78 2194 82
rect 2438 78 2442 82
rect 2526 78 2530 82
rect 2614 78 2618 82
rect 2734 78 2738 82
rect 2870 78 2874 82
rect 2990 78 2994 82
rect 2998 78 3002 82
rect 3078 78 3082 82
rect 3214 78 3218 82
rect 3430 78 3434 82
rect 3606 78 3610 82
rect 3630 78 3634 82
rect 3710 78 3714 82
rect 3806 78 3810 82
rect 4166 78 4170 82
rect 30 68 34 72
rect 158 68 162 72
rect 254 68 258 72
rect 542 68 546 72
rect 638 68 642 72
rect 734 68 738 72
rect 870 68 874 72
rect 918 68 922 72
rect 998 68 1002 72
rect 1014 68 1018 72
rect 1030 68 1034 72
rect 1102 68 1106 72
rect 1126 68 1130 72
rect 1214 68 1218 72
rect 1311 68 1315 72
rect 1326 68 1330 72
rect 1374 68 1378 72
rect 1398 68 1402 72
rect 1502 68 1506 72
rect 1662 68 1666 72
rect 1718 68 1722 72
rect 1894 68 1898 72
rect 1982 68 1986 72
rect 2054 68 2058 72
rect 2062 68 2066 72
rect 2150 68 2154 72
rect 2158 68 2162 72
rect 2238 68 2242 72
rect 2326 68 2330 72
rect 2414 68 2418 72
rect 2542 68 2546 72
rect 2630 68 2634 72
rect 2670 68 2674 72
rect 2678 68 2682 72
rect 2758 68 2762 72
rect 2774 68 2778 72
rect 2886 68 2890 72
rect 2974 68 2978 72
rect 3038 68 3042 72
rect 3094 68 3098 72
rect 3166 68 3170 72
rect 3206 68 3210 72
rect 3222 68 3226 72
rect 3238 68 3242 72
rect 3254 68 3258 72
rect 3334 68 3338 72
rect 3446 68 3450 72
rect 3534 68 3538 72
rect 3638 68 3642 72
rect 3678 68 3682 72
rect 3694 68 3698 72
rect 3725 68 3729 72
rect 3822 68 3826 72
rect 3958 68 3962 72
rect 3966 68 3970 72
rect 4118 68 4122 72
rect 4142 68 4146 72
rect 4198 68 4202 72
rect 4206 68 4210 72
rect 22 58 26 62
rect 198 58 202 62
rect 230 58 234 62
rect 342 58 346 62
rect 350 58 354 62
rect 374 58 378 62
rect 414 58 418 62
rect 445 58 449 62
rect 582 58 586 62
rect 630 58 634 62
rect 638 58 642 62
rect 686 58 690 62
rect 862 58 866 62
rect 878 58 882 62
rect 926 58 930 62
rect 974 58 978 62
rect 1006 58 1010 62
rect 1038 58 1042 62
rect 1086 58 1090 62
rect 1166 58 1170 62
rect 1366 58 1370 62
rect 1558 58 1562 62
rect 1766 58 1770 62
rect 1838 58 1842 62
rect 1966 58 1970 62
rect 2006 58 2010 62
rect 2014 58 2018 62
rect 2030 58 2034 62
rect 2206 58 2210 62
rect 2214 58 2218 62
rect 2270 58 2274 62
rect 2302 58 2306 62
rect 2334 58 2338 62
rect 2358 58 2362 62
rect 2486 58 2490 62
rect 2582 58 2586 62
rect 2622 58 2626 62
rect 2646 58 2650 62
rect 2662 58 2666 62
rect 2686 58 2690 62
rect 2710 58 2714 62
rect 2742 58 2746 62
rect 2774 58 2778 62
rect 2934 58 2938 62
rect 3142 58 3146 62
rect 3174 58 3178 62
rect 3190 58 3194 62
rect 3198 58 3202 62
rect 3230 58 3234 62
rect 3246 58 3250 62
rect 3502 58 3506 62
rect 3550 58 3554 62
rect 3558 58 3562 62
rect 3582 58 3586 62
rect 3614 58 3618 62
rect 3646 58 3650 62
rect 3670 58 3674 62
rect 3686 58 3690 62
rect 3766 58 3770 62
rect 3878 58 3882 62
rect 4054 58 4058 62
rect 4102 58 4106 62
rect 4134 58 4138 62
rect 4150 58 4154 62
rect 4190 58 4194 62
rect 4246 58 4250 62
rect 4278 58 4282 62
rect 4318 58 4322 62
rect 4342 58 4346 62
rect 190 50 194 54
rect 574 50 578 54
rect 614 48 618 52
rect 630 48 634 52
rect 702 50 706 54
rect 846 48 850 52
rect 862 48 866 52
rect 942 48 946 52
rect 1022 48 1026 52
rect 1054 48 1058 52
rect 1110 48 1114 52
rect 1182 50 1186 54
rect 1470 50 1474 54
rect 1750 50 1754 54
rect 1942 48 1946 52
rect 2006 48 2010 52
rect 2038 48 2042 52
rect 2134 48 2138 52
rect 2174 48 2178 52
rect 2310 48 2314 52
rect 2398 48 2402 52
rect 2574 50 2578 54
rect 2646 48 2650 52
rect 2662 48 2666 52
rect 2702 48 2706 52
rect 2934 48 2938 52
rect 3126 50 3130 54
rect 3190 48 3194 52
rect 3262 48 3266 52
rect 3494 48 3498 52
rect 3574 48 3578 52
rect 3606 48 3610 52
rect 3654 48 3658 52
rect 3670 48 3674 52
rect 3854 50 3858 54
rect 4166 48 4170 52
rect 4174 48 4178 52
rect 4310 48 4314 52
rect 6 38 10 42
rect 1086 38 1090 42
rect 1342 38 1346 42
rect 1398 38 1402 42
rect 1430 38 1434 42
rect 2150 38 2154 42
rect 4326 38 4330 42
rect 574 27 578 31
rect 702 27 706 31
rect 1182 27 1186 31
rect 1470 27 1474 31
rect 1750 27 1754 31
rect 3126 27 3130 31
rect 190 18 194 22
rect 246 18 250 22
rect 326 18 330 22
rect 366 18 370 22
rect 406 18 410 22
rect 430 18 434 22
rect 662 18 666 22
rect 894 18 898 22
rect 966 18 970 22
rect 990 18 994 22
rect 1078 18 1082 22
rect 1350 18 1354 22
rect 1942 18 1946 22
rect 2574 18 2578 22
rect 2934 18 2938 22
rect 3494 18 3498 22
rect 3854 18 3858 22
rect 4070 18 4074 22
rect 394 3 398 7
rect 401 3 405 7
rect 1418 3 1422 7
rect 1425 3 1429 7
rect 2442 3 2446 7
rect 2449 3 2453 7
rect 3474 3 3478 7
rect 3481 3 3485 7
<< metal2 >>
rect 1134 3128 1138 3132
rect 1158 3128 1162 3132
rect 1254 3128 1258 3132
rect 1358 3128 1362 3132
rect 1470 3128 1474 3132
rect 1558 3131 1562 3132
rect 1558 3128 1569 3131
rect 1638 3128 1642 3132
rect 1694 3128 1698 3132
rect 1726 3131 1730 3132
rect 1750 3131 1754 3132
rect 1774 3131 1778 3132
rect 1726 3128 1737 3131
rect 1750 3128 1761 3131
rect 896 3103 898 3107
rect 902 3103 905 3107
rect 909 3103 912 3107
rect 1134 3102 1137 3128
rect 1158 3102 1161 3128
rect 1254 3102 1257 3128
rect 1358 3102 1361 3128
rect 1470 3102 1473 3128
rect 650 3088 654 3091
rect 690 3088 694 3091
rect 618 3078 622 3081
rect 630 3078 638 3081
rect 642 3078 654 3081
rect 214 3072 217 3078
rect 230 3072 233 3078
rect 438 3072 441 3078
rect 454 3072 457 3078
rect 566 3072 569 3078
rect 74 3068 78 3071
rect 554 3068 558 3071
rect 6 3022 9 3068
rect 78 3062 81 3068
rect 230 3062 233 3068
rect 598 3062 601 3078
rect 610 3068 614 3071
rect 315 3058 318 3061
rect 562 3058 566 3061
rect 618 3058 622 3061
rect 6 2862 9 2928
rect 6 2762 9 2858
rect 14 2782 17 2818
rect 22 2781 25 2878
rect 30 2872 33 3058
rect 134 3002 137 3018
rect 110 2952 113 2978
rect 158 2962 161 3048
rect 182 3042 185 3050
rect 214 2960 217 3048
rect 270 3031 273 3058
rect 246 2952 249 2978
rect 62 2792 65 2908
rect 94 2842 97 2928
rect 110 2912 113 2938
rect 174 2882 177 2938
rect 246 2911 249 2938
rect 238 2908 249 2911
rect 262 2932 265 2998
rect 102 2872 105 2878
rect 158 2822 161 2828
rect 22 2778 33 2781
rect 22 2762 25 2768
rect 30 2752 33 2778
rect 38 2752 41 2758
rect 70 2752 73 2778
rect 86 2772 89 2818
rect 174 2782 177 2878
rect 238 2872 241 2908
rect 262 2902 265 2928
rect 274 2878 278 2881
rect 194 2868 201 2871
rect 198 2792 201 2868
rect 234 2858 238 2861
rect 214 2832 217 2848
rect 246 2832 249 2858
rect 254 2812 257 2868
rect 266 2858 270 2861
rect 310 2854 313 3048
rect 334 3042 337 3048
rect 350 2992 353 3058
rect 386 3048 390 3051
rect 494 3031 497 3058
rect 582 3052 585 3058
rect 538 3028 542 3031
rect 392 3003 394 3007
rect 398 3003 401 3007
rect 405 3003 408 3007
rect 478 2952 481 2988
rect 342 2948 343 2951
rect 347 2948 350 2951
rect 434 2948 438 2951
rect 342 2882 345 2948
rect 374 2942 377 2948
rect 354 2938 358 2941
rect 382 2932 385 2948
rect 542 2942 545 2948
rect 442 2928 446 2931
rect 414 2922 417 2928
rect 358 2882 361 2898
rect 302 2762 305 2828
rect 102 2752 105 2758
rect 158 2752 161 2758
rect 34 2738 38 2741
rect 50 2738 54 2741
rect 90 2738 94 2741
rect 146 2738 150 2741
rect 78 2732 81 2738
rect 102 2732 105 2738
rect 166 2732 169 2748
rect 62 2702 65 2728
rect 94 2712 97 2728
rect 118 2722 121 2728
rect 174 2722 177 2738
rect 182 2682 185 2728
rect 70 2672 73 2678
rect 38 2602 41 2650
rect 86 2622 89 2678
rect 190 2672 193 2758
rect 250 2738 254 2741
rect 222 2722 225 2728
rect 198 2692 201 2708
rect 126 2631 129 2658
rect 6 2542 9 2548
rect 22 2532 25 2548
rect 30 2542 33 2568
rect 94 2552 97 2588
rect 114 2558 118 2561
rect 118 2542 121 2548
rect 142 2542 145 2668
rect 198 2662 201 2688
rect 170 2648 174 2651
rect 206 2562 209 2708
rect 218 2678 222 2681
rect 230 2672 233 2688
rect 238 2672 241 2738
rect 270 2732 273 2748
rect 286 2742 289 2748
rect 278 2732 281 2738
rect 302 2712 305 2758
rect 314 2748 318 2751
rect 314 2738 318 2741
rect 326 2722 329 2788
rect 342 2772 345 2868
rect 398 2831 401 2858
rect 326 2692 329 2718
rect 214 2662 217 2668
rect 262 2662 265 2678
rect 318 2672 321 2678
rect 350 2672 353 2808
rect 392 2803 394 2807
rect 398 2803 401 2807
rect 405 2803 408 2807
rect 422 2792 425 2928
rect 558 2922 561 2938
rect 570 2928 574 2931
rect 430 2892 433 2918
rect 470 2872 473 2918
rect 478 2862 481 2868
rect 494 2861 497 2918
rect 518 2872 521 2898
rect 486 2858 497 2861
rect 502 2862 505 2868
rect 542 2862 545 2898
rect 550 2872 553 2918
rect 558 2882 561 2918
rect 566 2902 569 2918
rect 570 2878 574 2881
rect 582 2871 585 3048
rect 630 3032 633 3078
rect 678 3072 681 3088
rect 718 3072 721 3078
rect 798 3072 801 3078
rect 786 3068 790 3071
rect 654 3062 657 3068
rect 590 2952 593 2978
rect 622 2962 625 2978
rect 618 2948 622 2951
rect 606 2942 609 2948
rect 622 2932 625 2938
rect 630 2932 633 3028
rect 670 2952 673 3058
rect 694 3052 697 3058
rect 686 2952 689 2968
rect 682 2948 685 2951
rect 654 2942 657 2948
rect 670 2942 673 2948
rect 650 2928 654 2931
rect 646 2912 649 2928
rect 602 2878 606 2881
rect 634 2878 641 2881
rect 574 2868 585 2871
rect 438 2812 441 2818
rect 358 2672 361 2778
rect 430 2752 433 2778
rect 462 2762 465 2788
rect 430 2732 433 2738
rect 414 2722 417 2728
rect 386 2678 390 2681
rect 338 2668 342 2671
rect 250 2658 254 2661
rect 238 2632 241 2658
rect 250 2648 254 2651
rect 214 2572 217 2628
rect 262 2592 265 2658
rect 278 2652 281 2658
rect 274 2588 278 2591
rect 198 2552 201 2558
rect 206 2552 209 2558
rect 214 2552 217 2568
rect 234 2558 238 2561
rect 250 2548 254 2551
rect 190 2542 193 2548
rect 82 2538 86 2541
rect 154 2538 158 2541
rect 178 2538 182 2541
rect 266 2538 270 2541
rect 22 2352 25 2528
rect 110 2502 113 2518
rect 126 2502 129 2538
rect 214 2532 217 2538
rect 174 2502 177 2528
rect 230 2512 233 2528
rect 70 2472 73 2498
rect 166 2492 169 2498
rect 214 2492 217 2498
rect 86 2482 89 2488
rect 190 2482 193 2488
rect 238 2472 241 2518
rect 294 2492 297 2668
rect 358 2662 361 2668
rect 374 2662 377 2668
rect 414 2662 417 2708
rect 422 2692 425 2698
rect 442 2678 446 2681
rect 302 2652 305 2658
rect 414 2642 417 2658
rect 392 2603 394 2607
rect 398 2603 401 2607
rect 405 2603 408 2607
rect 374 2552 377 2578
rect 422 2562 425 2608
rect 358 2502 361 2528
rect 374 2482 377 2538
rect 390 2492 393 2508
rect 382 2482 385 2488
rect 294 2462 297 2478
rect 310 2472 313 2478
rect 410 2458 414 2461
rect 34 2450 38 2453
rect 126 2431 129 2458
rect 254 2431 257 2458
rect 362 2448 366 2451
rect 414 2442 417 2458
rect 422 2452 425 2558
rect 430 2532 433 2678
rect 454 2512 457 2668
rect 462 2662 465 2758
rect 470 2562 473 2818
rect 478 2762 481 2818
rect 486 2762 489 2858
rect 478 2692 481 2758
rect 486 2612 489 2758
rect 486 2592 489 2598
rect 470 2471 473 2558
rect 494 2542 497 2848
rect 502 2802 505 2848
rect 526 2792 529 2818
rect 534 2802 537 2838
rect 550 2782 553 2868
rect 558 2792 561 2858
rect 574 2852 577 2868
rect 590 2862 593 2868
rect 622 2862 625 2868
rect 574 2842 577 2848
rect 534 2762 537 2768
rect 502 2752 505 2758
rect 526 2752 529 2758
rect 506 2738 510 2741
rect 530 2738 534 2741
rect 518 2732 521 2738
rect 534 2692 537 2728
rect 550 2702 553 2758
rect 574 2752 577 2838
rect 582 2792 585 2858
rect 630 2842 633 2848
rect 590 2761 593 2818
rect 590 2758 598 2761
rect 574 2732 577 2738
rect 566 2722 569 2728
rect 558 2672 561 2708
rect 566 2692 569 2698
rect 506 2658 510 2661
rect 526 2652 529 2658
rect 526 2642 529 2648
rect 534 2642 537 2648
rect 510 2582 513 2618
rect 542 2592 545 2608
rect 550 2602 553 2658
rect 558 2652 561 2668
rect 582 2662 585 2748
rect 606 2742 609 2818
rect 578 2658 582 2661
rect 590 2652 593 2658
rect 570 2648 577 2651
rect 566 2592 569 2638
rect 514 2568 518 2571
rect 530 2568 534 2571
rect 518 2542 521 2548
rect 542 2542 545 2548
rect 490 2538 494 2541
rect 478 2501 481 2538
rect 498 2528 502 2531
rect 486 2512 489 2518
rect 550 2512 553 2558
rect 574 2532 577 2648
rect 590 2572 593 2648
rect 598 2582 601 2668
rect 606 2592 609 2728
rect 630 2692 633 2758
rect 638 2752 641 2878
rect 646 2872 649 2888
rect 654 2872 657 2918
rect 662 2872 665 2918
rect 670 2902 673 2938
rect 662 2862 665 2868
rect 694 2802 697 3048
rect 702 3032 705 3068
rect 734 3062 737 3068
rect 710 3052 713 3058
rect 790 3052 793 3068
rect 814 3062 817 3078
rect 838 3072 841 3088
rect 950 3072 953 3078
rect 882 3068 889 3071
rect 878 3062 881 3068
rect 842 3058 846 3061
rect 830 3052 833 3058
rect 858 3048 862 3051
rect 726 3042 729 3048
rect 750 3042 753 3048
rect 822 2982 825 3018
rect 782 2952 785 2978
rect 866 2958 870 2961
rect 830 2942 833 2958
rect 878 2952 881 2968
rect 766 2932 769 2938
rect 782 2932 785 2938
rect 710 2831 713 2858
rect 742 2792 745 2818
rect 686 2772 689 2778
rect 674 2758 678 2761
rect 722 2758 726 2761
rect 750 2752 753 2878
rect 766 2862 769 2868
rect 814 2852 817 2938
rect 854 2912 857 2928
rect 838 2892 841 2898
rect 870 2892 873 2948
rect 886 2942 889 3068
rect 926 3032 929 3058
rect 954 3048 958 3051
rect 942 3042 945 3048
rect 926 2942 929 3028
rect 974 2962 977 2968
rect 902 2922 905 2928
rect 926 2912 929 2938
rect 942 2932 945 2938
rect 950 2932 953 2958
rect 974 2942 977 2958
rect 958 2922 961 2938
rect 974 2912 977 2918
rect 896 2903 898 2907
rect 902 2903 905 2907
rect 909 2903 912 2907
rect 926 2892 929 2898
rect 758 2752 761 2758
rect 806 2752 809 2798
rect 738 2748 742 2751
rect 718 2732 721 2748
rect 742 2742 745 2748
rect 798 2742 801 2748
rect 698 2728 702 2731
rect 618 2648 622 2651
rect 614 2632 617 2648
rect 638 2612 641 2658
rect 646 2592 649 2648
rect 662 2622 665 2718
rect 750 2712 753 2738
rect 782 2732 785 2738
rect 806 2732 809 2748
rect 774 2722 777 2728
rect 594 2548 598 2551
rect 562 2528 566 2531
rect 478 2498 489 2501
rect 486 2492 489 2498
rect 470 2468 478 2471
rect 392 2403 394 2407
rect 398 2403 401 2407
rect 405 2403 408 2407
rect 438 2392 441 2418
rect 182 2362 185 2388
rect 310 2360 313 2379
rect 186 2348 190 2351
rect 290 2348 294 2351
rect 6 2292 9 2348
rect 134 2342 137 2348
rect 26 2338 30 2341
rect 210 2338 214 2341
rect 118 2322 121 2328
rect 22 2272 25 2308
rect 62 2282 65 2288
rect 174 2282 177 2288
rect 190 2272 193 2288
rect 26 2268 30 2271
rect 38 2262 41 2268
rect 222 2262 225 2348
rect 342 2332 345 2338
rect 358 2332 361 2358
rect 470 2342 473 2468
rect 478 2392 481 2428
rect 494 2412 497 2478
rect 502 2472 505 2478
rect 542 2462 545 2508
rect 566 2492 569 2508
rect 574 2492 577 2528
rect 582 2482 585 2528
rect 590 2492 593 2538
rect 606 2492 609 2508
rect 622 2492 625 2548
rect 586 2478 590 2481
rect 550 2472 553 2478
rect 506 2448 510 2451
rect 526 2422 529 2448
rect 558 2412 561 2478
rect 630 2472 633 2568
rect 642 2528 646 2531
rect 642 2488 646 2491
rect 618 2458 622 2461
rect 574 2422 577 2458
rect 610 2448 614 2451
rect 518 2360 521 2379
rect 610 2348 614 2351
rect 262 2282 265 2318
rect 358 2301 361 2328
rect 350 2298 361 2301
rect 350 2282 353 2298
rect 6 2252 9 2258
rect 22 2252 25 2258
rect 38 2242 41 2248
rect 54 2222 57 2228
rect 54 2182 57 2188
rect 6 2172 9 2178
rect 30 2162 33 2168
rect 70 2152 73 2158
rect 222 2152 225 2258
rect 238 2222 241 2248
rect 366 2242 369 2268
rect 418 2258 422 2261
rect 398 2222 401 2250
rect 270 2192 273 2218
rect 392 2203 394 2207
rect 398 2203 401 2207
rect 405 2203 408 2207
rect 230 2162 233 2188
rect 254 2162 257 2188
rect 310 2162 313 2168
rect 262 2152 265 2158
rect 26 2148 30 2151
rect 50 2148 54 2151
rect 82 2148 85 2151
rect 306 2148 310 2151
rect 182 2142 185 2148
rect 166 2132 169 2138
rect 30 2052 33 2068
rect 46 2062 49 2118
rect 166 2082 169 2088
rect 182 2072 185 2098
rect 82 2068 85 2071
rect 54 2052 57 2068
rect 62 2062 65 2068
rect 230 2062 233 2148
rect 286 2082 289 2138
rect 294 2122 297 2148
rect 318 2142 321 2188
rect 366 2162 369 2188
rect 338 2148 342 2151
rect 334 2092 337 2128
rect 334 2082 337 2088
rect 318 2062 321 2068
rect 374 2062 377 2148
rect 414 2112 417 2138
rect 430 2132 433 2338
rect 462 2252 465 2258
rect 430 2082 433 2128
rect 470 2092 473 2328
rect 550 2312 553 2338
rect 566 2332 569 2338
rect 566 2302 569 2328
rect 534 2282 537 2298
rect 606 2272 609 2348
rect 622 2272 625 2418
rect 646 2392 649 2478
rect 654 2472 657 2528
rect 662 2332 665 2618
rect 670 2592 673 2658
rect 678 2654 681 2698
rect 806 2692 809 2718
rect 814 2702 817 2848
rect 838 2762 841 2848
rect 854 2842 857 2868
rect 874 2858 878 2861
rect 898 2858 902 2861
rect 822 2752 825 2758
rect 854 2752 857 2838
rect 870 2812 873 2848
rect 870 2772 873 2808
rect 862 2752 865 2768
rect 830 2742 833 2748
rect 870 2742 873 2748
rect 854 2732 857 2738
rect 834 2728 838 2731
rect 846 2701 849 2718
rect 838 2698 849 2701
rect 710 2672 713 2678
rect 726 2662 729 2678
rect 814 2672 817 2678
rect 838 2662 841 2698
rect 854 2692 857 2708
rect 846 2682 849 2688
rect 846 2672 849 2678
rect 854 2672 857 2688
rect 862 2662 865 2738
rect 870 2722 873 2728
rect 878 2692 881 2848
rect 910 2752 913 2758
rect 918 2752 921 2878
rect 942 2862 945 2888
rect 950 2872 953 2908
rect 982 2892 985 3038
rect 998 3031 1001 3058
rect 1038 3032 1041 3078
rect 1054 3072 1057 3078
rect 1198 3072 1201 3098
rect 1270 3072 1273 3098
rect 1290 3058 1294 3061
rect 1106 3048 1110 3051
rect 1134 3042 1137 3048
rect 1150 2992 1153 3058
rect 1174 3042 1177 3058
rect 1266 3038 1270 3041
rect 994 2958 998 2961
rect 1030 2952 1033 2988
rect 1142 2952 1145 2978
rect 1174 2962 1177 3038
rect 1294 3022 1297 3048
rect 1182 2992 1185 3018
rect 1002 2948 1006 2951
rect 1002 2938 1006 2941
rect 1010 2888 1014 2891
rect 1038 2882 1041 2928
rect 1046 2892 1049 2928
rect 1038 2872 1041 2878
rect 962 2868 966 2871
rect 926 2842 929 2848
rect 950 2821 953 2868
rect 942 2818 953 2821
rect 886 2722 889 2748
rect 894 2742 897 2748
rect 906 2728 910 2731
rect 766 2631 769 2658
rect 822 2592 825 2648
rect 854 2592 857 2648
rect 790 2582 793 2588
rect 810 2558 817 2561
rect 834 2558 838 2561
rect 726 2542 729 2548
rect 670 2362 673 2518
rect 790 2502 793 2518
rect 814 2492 817 2558
rect 862 2552 865 2658
rect 826 2548 830 2551
rect 870 2542 873 2688
rect 886 2682 889 2718
rect 896 2703 898 2707
rect 902 2703 905 2707
rect 909 2703 912 2707
rect 898 2688 902 2691
rect 942 2682 945 2818
rect 950 2732 953 2768
rect 966 2742 969 2858
rect 982 2842 985 2848
rect 990 2772 993 2868
rect 1062 2862 1065 2878
rect 1078 2872 1081 2908
rect 1070 2862 1073 2868
rect 1058 2858 1062 2861
rect 974 2742 977 2748
rect 982 2732 985 2738
rect 990 2722 993 2758
rect 1002 2748 1006 2751
rect 1014 2742 1017 2768
rect 1046 2752 1049 2848
rect 1042 2748 1046 2751
rect 1022 2742 1025 2748
rect 1054 2742 1057 2748
rect 1002 2738 1006 2741
rect 1022 2722 1025 2728
rect 950 2682 953 2718
rect 942 2672 945 2678
rect 922 2668 926 2671
rect 958 2661 961 2718
rect 1046 2712 1049 2718
rect 954 2658 961 2661
rect 898 2648 902 2651
rect 878 2602 881 2648
rect 998 2631 1001 2658
rect 918 2560 921 2579
rect 950 2542 953 2548
rect 834 2538 838 2541
rect 966 2532 969 2568
rect 896 2503 898 2507
rect 902 2503 905 2507
rect 909 2503 912 2507
rect 726 2442 729 2478
rect 814 2472 817 2488
rect 926 2482 929 2488
rect 1006 2482 1009 2548
rect 1038 2502 1041 2678
rect 1054 2672 1057 2678
rect 1086 2654 1089 2938
rect 1126 2842 1129 2928
rect 1142 2902 1145 2938
rect 1206 2872 1209 3018
rect 1230 2962 1233 2988
rect 1342 2982 1345 3068
rect 1238 2952 1241 2958
rect 1278 2932 1281 2938
rect 1294 2922 1297 2928
rect 1358 2902 1361 3078
rect 1538 3068 1542 3071
rect 1398 2992 1401 3058
rect 1534 3022 1537 3068
rect 1558 3022 1561 3048
rect 1416 3003 1418 3007
rect 1422 3003 1425 3007
rect 1429 3003 1432 3007
rect 1410 2948 1414 2951
rect 1390 2932 1393 2938
rect 1270 2882 1273 2898
rect 1126 2802 1129 2818
rect 1182 2812 1185 2868
rect 1254 2862 1257 2868
rect 1150 2792 1153 2798
rect 1150 2732 1153 2788
rect 1166 2732 1169 2738
rect 1142 2692 1145 2708
rect 1150 2662 1153 2698
rect 1166 2692 1169 2718
rect 1182 2692 1185 2708
rect 1198 2662 1201 2828
rect 1206 2752 1209 2858
rect 1222 2831 1225 2850
rect 1214 2762 1217 2788
rect 1206 2722 1209 2748
rect 1214 2692 1217 2728
rect 1210 2668 1214 2671
rect 1046 2592 1049 2598
rect 742 2462 745 2468
rect 726 2422 729 2438
rect 774 2431 777 2450
rect 782 2352 785 2458
rect 878 2431 881 2450
rect 814 2360 817 2379
rect 726 2342 729 2348
rect 766 2332 769 2338
rect 690 2318 694 2321
rect 662 2272 665 2318
rect 670 2282 673 2318
rect 650 2268 654 2271
rect 518 2262 521 2268
rect 574 2262 577 2268
rect 670 2262 673 2278
rect 694 2272 697 2308
rect 710 2272 713 2318
rect 682 2268 686 2271
rect 730 2268 734 2271
rect 486 2231 489 2250
rect 510 2192 513 2218
rect 537 2138 545 2141
rect 530 2128 537 2131
rect 518 2092 521 2108
rect 234 2058 238 2061
rect 266 2058 270 2061
rect 6 2042 9 2048
rect 6 1992 9 2008
rect 70 1992 73 2018
rect 34 1988 38 1991
rect 62 1962 65 1968
rect 78 1962 81 1968
rect 22 1952 25 1958
rect 50 1948 54 1951
rect 66 1948 70 1951
rect 86 1942 89 2048
rect 214 2022 217 2050
rect 142 1992 145 1998
rect 122 1978 126 1981
rect 222 1962 225 1978
rect 98 1958 102 1961
rect 178 1958 182 1961
rect 98 1948 102 1951
rect 54 1882 57 1938
rect 86 1932 89 1938
rect 30 1872 33 1878
rect 54 1872 57 1878
rect 62 1862 65 1898
rect 86 1882 89 1928
rect 110 1892 113 1958
rect 134 1952 137 1958
rect 158 1942 161 1948
rect 174 1942 177 1948
rect 166 1932 169 1938
rect 190 1922 193 1958
rect 206 1952 209 1958
rect 230 1952 233 1968
rect 238 1962 241 1968
rect 198 1932 201 1938
rect 206 1902 209 1948
rect 230 1942 233 1948
rect 218 1938 222 1941
rect 26 1858 30 1861
rect 74 1858 78 1861
rect 54 1852 57 1858
rect 90 1848 94 1851
rect 6 1842 9 1848
rect 78 1832 81 1848
rect 30 1772 33 1778
rect 22 1752 25 1758
rect 6 1742 9 1748
rect 34 1688 38 1691
rect 6 1672 9 1678
rect 26 1658 30 1661
rect 102 1592 105 1878
rect 174 1852 177 1878
rect 190 1872 193 1878
rect 246 1862 249 2058
rect 286 2031 289 2050
rect 392 2003 394 2007
rect 398 2003 401 2007
rect 405 2003 408 2007
rect 253 1942 256 1948
rect 350 1942 353 1968
rect 398 1962 401 1988
rect 334 1932 337 1938
rect 262 1872 265 1918
rect 290 1888 294 1891
rect 366 1882 369 1908
rect 398 1902 401 1948
rect 422 1892 425 2078
rect 446 2072 449 2088
rect 534 2072 537 2128
rect 542 2112 545 2138
rect 550 2092 553 2198
rect 574 2152 577 2258
rect 670 2222 673 2248
rect 614 2192 617 2218
rect 638 2212 641 2218
rect 614 2142 617 2178
rect 678 2162 681 2188
rect 614 2132 617 2138
rect 630 2132 633 2138
rect 606 2072 609 2078
rect 614 2072 617 2108
rect 646 2082 649 2088
rect 654 2072 657 2108
rect 678 2092 681 2138
rect 686 2112 689 2268
rect 722 2258 726 2261
rect 742 2261 745 2298
rect 750 2292 753 2308
rect 782 2292 785 2338
rect 822 2302 825 2418
rect 910 2402 913 2468
rect 966 2462 969 2478
rect 834 2348 838 2351
rect 822 2272 825 2278
rect 762 2268 766 2271
rect 738 2258 745 2261
rect 762 2258 766 2261
rect 810 2258 814 2261
rect 826 2258 830 2261
rect 842 2258 846 2261
rect 706 2248 710 2251
rect 818 2248 822 2251
rect 750 2192 753 2248
rect 774 2192 777 2228
rect 782 2211 785 2248
rect 790 2242 793 2248
rect 846 2242 849 2248
rect 862 2242 865 2368
rect 878 2352 881 2358
rect 886 2292 889 2398
rect 902 2360 905 2379
rect 990 2352 993 2478
rect 1046 2472 1049 2478
rect 1006 2468 1007 2471
rect 1011 2468 1014 2472
rect 934 2332 937 2338
rect 950 2311 953 2328
rect 942 2308 953 2311
rect 896 2303 898 2307
rect 902 2303 905 2307
rect 909 2303 912 2307
rect 902 2262 905 2278
rect 914 2268 918 2271
rect 926 2262 929 2268
rect 874 2258 878 2261
rect 934 2252 937 2298
rect 798 2232 801 2238
rect 862 2232 865 2238
rect 782 2208 809 2211
rect 806 2192 809 2208
rect 710 2161 713 2188
rect 742 2172 745 2178
rect 814 2172 817 2178
rect 722 2168 726 2171
rect 710 2158 721 2161
rect 702 2152 705 2158
rect 686 2092 689 2098
rect 710 2072 713 2138
rect 718 2072 721 2158
rect 726 2082 729 2088
rect 466 2068 470 2071
rect 498 2068 502 2071
rect 482 2058 486 2061
rect 506 2058 510 2061
rect 522 2058 526 2061
rect 626 2058 630 2061
rect 446 1942 449 1978
rect 449 1938 454 1941
rect 382 1872 385 1878
rect 190 1752 193 1858
rect 238 1822 241 1848
rect 262 1792 265 1868
rect 278 1842 281 1848
rect 242 1788 246 1791
rect 206 1762 209 1788
rect 158 1742 161 1748
rect 142 1732 145 1738
rect 142 1642 145 1678
rect 158 1672 161 1678
rect 206 1662 209 1748
rect 334 1742 337 1768
rect 366 1760 369 1779
rect 382 1752 385 1858
rect 414 1822 417 1850
rect 392 1803 394 1807
rect 398 1803 401 1807
rect 405 1803 408 1807
rect 422 1742 425 1888
rect 430 1862 433 1898
rect 434 1858 438 1861
rect 462 1792 465 1828
rect 470 1822 473 2058
rect 662 2052 665 2058
rect 522 2048 526 2051
rect 626 2048 630 2051
rect 486 2042 489 2048
rect 678 2032 681 2048
rect 630 2012 633 2018
rect 622 1992 625 1998
rect 574 1960 577 1979
rect 638 1972 641 1978
rect 654 1962 657 1968
rect 638 1952 641 1958
rect 662 1952 665 1998
rect 686 1982 689 2048
rect 694 1992 697 1998
rect 702 1992 705 2058
rect 710 1972 713 2068
rect 734 2052 737 2168
rect 742 2052 745 2168
rect 758 2162 761 2168
rect 798 2162 801 2168
rect 770 2148 774 2151
rect 750 2132 753 2148
rect 790 2142 793 2158
rect 762 2138 766 2141
rect 766 2092 769 2128
rect 806 2112 809 2148
rect 814 2142 817 2168
rect 786 2068 790 2071
rect 754 2058 758 2061
rect 782 2052 785 2058
rect 770 2048 774 2051
rect 686 1962 689 1968
rect 682 1948 686 1951
rect 542 1942 545 1948
rect 526 1922 529 1928
rect 534 1872 537 1878
rect 550 1872 553 1878
rect 590 1862 593 1948
rect 614 1942 617 1948
rect 702 1942 705 1968
rect 710 1942 713 1948
rect 634 1938 638 1941
rect 658 1938 662 1941
rect 630 1892 633 1908
rect 638 1872 641 1938
rect 478 1852 481 1858
rect 486 1822 489 1848
rect 434 1758 438 1761
rect 450 1758 454 1761
rect 270 1692 273 1728
rect 318 1722 321 1728
rect 246 1662 249 1668
rect 210 1658 214 1661
rect 230 1652 233 1658
rect 206 1622 209 1648
rect 6 1582 9 1588
rect 30 1582 33 1588
rect 126 1572 129 1578
rect 234 1568 238 1571
rect 22 1552 25 1568
rect 142 1562 145 1568
rect 54 1558 62 1561
rect 82 1558 86 1561
rect 54 1552 57 1558
rect 66 1548 70 1551
rect 130 1548 134 1551
rect 6 1492 9 1498
rect 6 1422 9 1468
rect 30 1452 33 1478
rect 6 1372 9 1378
rect 22 1352 25 1358
rect 30 1352 33 1368
rect 18 1218 25 1221
rect 22 1152 25 1218
rect 38 1192 41 1498
rect 54 1472 57 1538
rect 62 1472 65 1478
rect 50 1468 54 1471
rect 70 1461 73 1548
rect 78 1502 81 1548
rect 146 1538 150 1541
rect 218 1538 222 1541
rect 166 1482 169 1518
rect 82 1478 86 1481
rect 182 1472 185 1478
rect 66 1458 73 1461
rect 78 1462 81 1468
rect 254 1462 257 1648
rect 270 1492 273 1548
rect 310 1542 313 1638
rect 318 1592 321 1718
rect 382 1672 385 1678
rect 338 1668 342 1671
rect 362 1668 366 1671
rect 326 1642 329 1668
rect 378 1658 382 1661
rect 326 1542 329 1578
rect 310 1532 313 1538
rect 358 1502 361 1658
rect 390 1652 393 1678
rect 422 1672 425 1738
rect 398 1642 401 1668
rect 430 1662 433 1748
rect 466 1718 470 1721
rect 486 1672 489 1718
rect 502 1682 505 1798
rect 590 1752 593 1858
rect 606 1762 609 1788
rect 610 1748 614 1751
rect 542 1732 545 1738
rect 478 1662 481 1668
rect 392 1603 394 1607
rect 398 1603 401 1607
rect 405 1603 408 1607
rect 422 1592 425 1598
rect 270 1482 273 1488
rect 366 1482 369 1588
rect 374 1562 377 1588
rect 382 1542 385 1548
rect 398 1542 401 1568
rect 430 1552 433 1658
rect 502 1642 505 1648
rect 478 1562 481 1588
rect 430 1542 433 1548
rect 302 1462 305 1478
rect 350 1472 353 1478
rect 46 1352 49 1368
rect 54 1352 57 1458
rect 182 1421 185 1458
rect 230 1422 233 1448
rect 182 1418 193 1421
rect 90 1388 94 1391
rect 62 1372 65 1378
rect 78 1362 81 1368
rect 102 1352 105 1378
rect 134 1362 137 1398
rect 146 1378 150 1381
rect 122 1358 126 1361
rect 114 1348 118 1351
rect 106 1338 110 1341
rect 54 1252 57 1338
rect 94 1272 97 1278
rect 110 1262 113 1268
rect 110 1192 113 1248
rect 142 1222 145 1250
rect 38 1172 41 1188
rect 86 1152 89 1158
rect 94 1152 97 1168
rect 126 1152 129 1198
rect 138 1148 142 1151
rect 62 1142 65 1148
rect 126 1122 129 1138
rect 150 1112 153 1158
rect 158 1152 161 1258
rect 182 1152 185 1388
rect 190 1352 193 1418
rect 254 1392 257 1458
rect 302 1422 305 1448
rect 294 1362 297 1388
rect 342 1382 345 1398
rect 346 1378 350 1381
rect 190 1262 193 1348
rect 230 1332 233 1358
rect 302 1352 305 1358
rect 246 1332 249 1338
rect 194 1258 198 1261
rect 198 1222 201 1248
rect 206 1162 209 1188
rect 202 1148 206 1151
rect 158 1142 161 1148
rect 182 1101 185 1148
rect 182 1098 190 1101
rect 6 1082 9 1088
rect 30 1072 33 1078
rect 142 1072 145 1078
rect 158 1072 161 1078
rect 6 1052 9 1068
rect 198 1062 201 1148
rect 26 1058 30 1061
rect 34 988 38 991
rect 6 972 9 978
rect 22 952 25 958
rect 198 952 201 1058
rect 206 1022 209 1048
rect 206 962 209 988
rect 158 942 161 948
rect 142 922 145 928
rect 142 882 145 888
rect 6 872 9 878
rect 30 862 33 868
rect 158 862 161 868
rect 22 852 25 858
rect 46 842 49 858
rect 58 848 62 851
rect 34 788 38 791
rect 6 772 9 778
rect 22 752 25 768
rect 198 752 201 858
rect 206 822 209 848
rect 206 762 209 788
rect 158 742 161 748
rect 142 722 145 728
rect 6 642 9 648
rect 118 632 121 678
rect 134 672 137 678
rect 78 542 81 548
rect 10 538 14 541
rect 6 442 9 448
rect 6 342 9 348
rect 14 342 17 538
rect 62 482 65 518
rect 118 482 121 618
rect 86 392 89 408
rect 26 348 30 351
rect 34 338 38 341
rect 18 218 25 221
rect 6 142 9 148
rect 22 62 25 218
rect 38 192 41 338
rect 94 282 97 388
rect 106 348 109 351
rect 118 322 121 478
rect 134 472 137 628
rect 150 562 153 608
rect 166 592 169 708
rect 198 672 201 748
rect 214 732 217 1298
rect 262 1282 265 1288
rect 358 1272 361 1388
rect 366 1362 369 1478
rect 454 1442 457 1548
rect 478 1542 481 1548
rect 526 1542 529 1588
rect 542 1532 545 1718
rect 558 1712 561 1738
rect 638 1692 641 1868
rect 654 1862 657 1878
rect 654 1842 657 1858
rect 646 1762 649 1788
rect 654 1782 657 1838
rect 662 1772 665 1858
rect 686 1852 689 1938
rect 710 1862 713 1868
rect 698 1858 702 1861
rect 718 1851 721 2048
rect 734 1991 737 2048
rect 742 2032 745 2038
rect 726 1988 737 1991
rect 726 1972 729 1988
rect 738 1978 742 1981
rect 750 1971 753 2038
rect 766 1992 769 1998
rect 774 1972 777 1978
rect 746 1968 753 1971
rect 790 1971 793 2068
rect 798 2052 801 2088
rect 810 2058 814 2061
rect 822 2042 825 2178
rect 838 2172 841 2178
rect 846 2172 849 2178
rect 862 2172 865 2228
rect 870 2192 873 2218
rect 878 2181 881 2248
rect 870 2178 881 2181
rect 830 2162 833 2168
rect 870 2161 873 2178
rect 866 2158 873 2161
rect 842 2148 846 2151
rect 838 2092 841 2138
rect 862 2092 865 2158
rect 870 2142 873 2148
rect 878 2132 881 2168
rect 934 2162 937 2248
rect 942 2202 945 2308
rect 958 2272 961 2278
rect 974 2272 977 2278
rect 982 2272 985 2308
rect 1006 2292 1009 2338
rect 1030 2332 1033 2418
rect 1054 2392 1057 2468
rect 1070 2462 1073 2608
rect 1126 2602 1129 2658
rect 1150 2612 1153 2658
rect 1182 2642 1185 2648
rect 1198 2602 1201 2658
rect 1210 2648 1214 2651
rect 1102 2552 1105 2558
rect 1094 2542 1097 2548
rect 1110 2542 1113 2588
rect 1122 2548 1126 2551
rect 1078 2522 1081 2538
rect 1222 2532 1225 2808
rect 1246 2792 1249 2808
rect 1270 2802 1273 2878
rect 1366 2862 1369 2868
rect 1374 2852 1377 2918
rect 1242 2668 1246 2671
rect 1254 2651 1257 2768
rect 1302 2760 1305 2779
rect 1350 2762 1353 2838
rect 1374 2832 1377 2838
rect 1382 2812 1385 2868
rect 1390 2782 1393 2928
rect 1398 2902 1401 2948
rect 1410 2938 1414 2941
rect 1426 2938 1430 2941
rect 1438 2922 1441 3018
rect 1478 2972 1481 3018
rect 1534 2972 1537 2978
rect 1462 2952 1465 2958
rect 1474 2948 1478 2951
rect 1410 2888 1414 2891
rect 1422 2882 1425 2918
rect 1430 2892 1433 2898
rect 1454 2892 1457 2948
rect 1470 2942 1473 2948
rect 1478 2932 1481 2938
rect 1486 2912 1489 2938
rect 1494 2932 1497 2948
rect 1494 2882 1497 2928
rect 1510 2922 1513 2958
rect 1534 2952 1537 2958
rect 1558 2942 1561 2978
rect 1538 2938 1542 2941
rect 1546 2928 1550 2931
rect 1558 2922 1561 2938
rect 1566 2892 1569 3128
rect 1694 3102 1697 3128
rect 1734 3092 1737 3128
rect 1758 3092 1761 3128
rect 1766 3128 1778 3131
rect 1798 3131 1802 3132
rect 1798 3128 1809 3131
rect 1766 3092 1769 3128
rect 1806 3092 1809 3128
rect 1902 3128 1906 3132
rect 1918 3128 1922 3132
rect 1998 3128 2002 3132
rect 2014 3131 2018 3132
rect 2038 3131 2042 3132
rect 2062 3131 2066 3132
rect 2014 3128 2025 3131
rect 2038 3128 2049 3131
rect 2062 3128 2073 3131
rect 1902 3102 1905 3128
rect 1918 3102 1921 3128
rect 1928 3103 1930 3107
rect 1934 3103 1937 3107
rect 1941 3103 1944 3107
rect 1894 3082 1897 3088
rect 1606 3062 1609 3068
rect 1582 2962 1585 2968
rect 1622 2942 1625 3078
rect 1878 3062 1881 3068
rect 1666 3058 1670 3061
rect 1630 2962 1633 2988
rect 1638 2952 1641 2988
rect 1678 2942 1681 2948
rect 1574 2932 1577 2938
rect 1582 2892 1585 2918
rect 1598 2912 1601 2938
rect 1606 2932 1609 2938
rect 1694 2932 1697 2938
rect 1638 2892 1641 2928
rect 1406 2852 1409 2878
rect 1438 2872 1441 2878
rect 1542 2872 1545 2888
rect 1638 2872 1641 2888
rect 1654 2862 1657 2908
rect 1466 2858 1470 2861
rect 1416 2803 1418 2807
rect 1422 2803 1425 2807
rect 1429 2803 1432 2807
rect 1446 2772 1449 2858
rect 1462 2792 1465 2848
rect 1486 2812 1489 2818
rect 1282 2748 1286 2751
rect 1262 2742 1265 2748
rect 1334 2732 1337 2738
rect 1350 2732 1353 2758
rect 1502 2752 1505 2828
rect 1542 2792 1545 2858
rect 1674 2848 1678 2851
rect 1666 2838 1670 2841
rect 1522 2788 1526 2791
rect 1646 2772 1649 2818
rect 1662 2762 1665 2788
rect 1686 2762 1689 2818
rect 1702 2792 1705 2908
rect 1742 2882 1745 3058
rect 1782 2992 1785 3058
rect 1790 2982 1793 3058
rect 1830 3022 1833 3048
rect 1798 2992 1801 2998
rect 1718 2792 1721 2878
rect 1750 2871 1753 2928
rect 1746 2868 1753 2871
rect 1774 2872 1777 2918
rect 1790 2882 1793 2978
rect 1814 2872 1817 2958
rect 1838 2952 1841 3058
rect 1942 2962 1945 2988
rect 1838 2902 1841 2948
rect 1878 2922 1881 2928
rect 1894 2912 1897 2938
rect 1966 2932 1969 2938
rect 1928 2903 1930 2907
rect 1934 2903 1937 2907
rect 1941 2903 1944 2907
rect 1814 2862 1817 2868
rect 1846 2862 1849 2868
rect 1886 2862 1889 2898
rect 1950 2882 1953 2888
rect 1934 2862 1937 2868
rect 1842 2858 1846 2861
rect 1750 2822 1753 2858
rect 1770 2848 1774 2851
rect 1670 2752 1673 2758
rect 1498 2748 1502 2751
rect 1250 2648 1257 2651
rect 1262 2672 1265 2688
rect 1334 2672 1337 2678
rect 1246 2592 1249 2648
rect 1262 2622 1265 2668
rect 1350 2662 1353 2678
rect 1390 2662 1393 2748
rect 1430 2692 1433 2718
rect 1270 2560 1273 2579
rect 1286 2552 1289 2658
rect 1302 2631 1305 2650
rect 1434 2618 1438 2621
rect 1238 2532 1241 2538
rect 1142 2522 1145 2528
rect 1150 2482 1153 2498
rect 1222 2492 1225 2528
rect 1086 2462 1089 2478
rect 1134 2462 1137 2468
rect 1066 2458 1070 2461
rect 1054 2342 1057 2348
rect 1030 2282 1033 2318
rect 1046 2312 1049 2338
rect 1062 2292 1065 2438
rect 1102 2431 1105 2450
rect 1126 2372 1129 2378
rect 1082 2368 1086 2371
rect 1042 2288 1046 2291
rect 950 2242 953 2258
rect 982 2241 985 2268
rect 982 2238 993 2241
rect 966 2222 969 2228
rect 954 2168 958 2171
rect 966 2162 969 2168
rect 922 2148 926 2151
rect 954 2148 958 2151
rect 906 2138 910 2141
rect 922 2138 926 2141
rect 938 2138 942 2141
rect 886 2092 889 2108
rect 896 2103 898 2107
rect 902 2103 905 2107
rect 909 2103 912 2107
rect 918 2092 921 2128
rect 974 2092 977 2118
rect 982 2092 985 2118
rect 942 2072 945 2078
rect 858 2068 862 2071
rect 810 2038 814 2041
rect 806 2022 809 2028
rect 830 1992 833 1998
rect 790 1968 801 1971
rect 726 1962 729 1968
rect 758 1962 761 1968
rect 734 1881 737 1948
rect 742 1892 745 1938
rect 766 1922 769 1948
rect 774 1891 777 1968
rect 790 1952 793 1958
rect 786 1918 790 1921
rect 766 1888 777 1891
rect 734 1878 745 1881
rect 726 1871 729 1878
rect 726 1868 734 1871
rect 730 1858 734 1861
rect 714 1848 721 1851
rect 702 1842 705 1848
rect 742 1842 745 1878
rect 766 1872 769 1888
rect 774 1872 777 1878
rect 798 1862 801 1968
rect 814 1952 817 1988
rect 838 1972 841 2018
rect 854 1992 857 2058
rect 862 2002 865 2068
rect 874 2058 878 2061
rect 886 2042 889 2048
rect 866 1978 870 1981
rect 822 1962 825 1968
rect 870 1952 873 1978
rect 878 1952 881 1988
rect 834 1948 838 1951
rect 806 1938 814 1941
rect 806 1902 809 1938
rect 806 1872 809 1898
rect 862 1882 865 1948
rect 918 1942 921 2068
rect 954 2058 958 2061
rect 934 1992 937 2058
rect 942 2022 945 2058
rect 966 2052 969 2078
rect 982 2062 985 2088
rect 990 2072 993 2238
rect 1006 2232 1009 2248
rect 1014 2192 1017 2278
rect 1054 2272 1057 2288
rect 1078 2262 1081 2358
rect 1094 2352 1097 2368
rect 1102 2352 1105 2358
rect 1086 2272 1089 2318
rect 1094 2292 1097 2328
rect 1110 2312 1113 2358
rect 1118 2272 1121 2358
rect 1134 2351 1137 2368
rect 1130 2348 1137 2351
rect 1034 2258 1038 2261
rect 1114 2258 1118 2261
rect 1078 2231 1081 2258
rect 1078 2228 1089 2231
rect 998 2152 1001 2158
rect 1014 2152 1017 2168
rect 1010 2138 1014 2141
rect 998 2072 1001 2088
rect 1006 2072 1009 2138
rect 926 1972 929 1978
rect 914 1938 918 1941
rect 886 1912 889 1938
rect 896 1903 898 1907
rect 902 1903 905 1907
rect 909 1903 912 1907
rect 826 1868 830 1871
rect 846 1862 849 1868
rect 854 1862 857 1878
rect 870 1871 873 1878
rect 886 1872 889 1898
rect 902 1872 905 1878
rect 926 1872 929 1948
rect 866 1868 873 1871
rect 918 1868 926 1871
rect 878 1862 881 1868
rect 918 1862 921 1868
rect 778 1858 782 1861
rect 758 1852 761 1858
rect 694 1772 697 1838
rect 742 1812 745 1818
rect 590 1672 593 1678
rect 606 1672 609 1678
rect 654 1662 657 1748
rect 694 1722 697 1738
rect 710 1732 713 1738
rect 702 1692 705 1708
rect 758 1692 761 1848
rect 782 1842 785 1848
rect 678 1672 681 1688
rect 606 1582 609 1658
rect 638 1622 641 1650
rect 582 1552 585 1578
rect 630 1542 633 1558
rect 638 1552 641 1598
rect 646 1572 649 1578
rect 662 1562 665 1618
rect 678 1562 681 1668
rect 718 1662 721 1668
rect 686 1642 689 1658
rect 714 1648 718 1651
rect 726 1642 729 1668
rect 742 1652 745 1688
rect 774 1672 777 1828
rect 798 1812 801 1848
rect 814 1822 817 1858
rect 794 1758 798 1761
rect 750 1652 753 1658
rect 694 1582 697 1588
rect 694 1552 697 1568
rect 670 1542 673 1548
rect 618 1538 623 1541
rect 690 1538 694 1541
rect 486 1482 489 1518
rect 486 1472 489 1478
rect 392 1403 394 1407
rect 398 1403 401 1407
rect 405 1403 408 1407
rect 378 1348 382 1351
rect 438 1342 441 1428
rect 470 1382 473 1468
rect 510 1462 513 1468
rect 518 1462 521 1478
rect 530 1468 534 1471
rect 498 1458 502 1461
rect 422 1302 425 1328
rect 478 1322 481 1458
rect 498 1448 502 1451
rect 534 1432 537 1438
rect 486 1362 489 1388
rect 526 1362 529 1388
rect 494 1352 497 1358
rect 522 1348 526 1351
rect 394 1268 398 1271
rect 246 1262 249 1268
rect 366 1232 369 1238
rect 374 1182 377 1268
rect 430 1262 433 1268
rect 462 1262 465 1308
rect 446 1252 449 1258
rect 454 1252 457 1258
rect 486 1252 489 1268
rect 498 1258 502 1261
rect 518 1252 521 1268
rect 526 1262 529 1268
rect 414 1212 417 1248
rect 534 1242 537 1398
rect 474 1238 478 1241
rect 506 1238 510 1241
rect 392 1203 394 1207
rect 398 1203 401 1207
rect 405 1203 408 1207
rect 454 1182 457 1218
rect 402 1178 406 1181
rect 354 1168 358 1171
rect 422 1162 425 1168
rect 430 1162 433 1168
rect 454 1152 457 1178
rect 462 1172 465 1218
rect 494 1161 497 1218
rect 490 1158 497 1161
rect 526 1161 529 1218
rect 522 1158 529 1161
rect 502 1152 505 1158
rect 534 1152 537 1158
rect 378 1148 382 1151
rect 442 1148 446 1151
rect 222 1071 225 1118
rect 254 1102 257 1138
rect 270 1122 273 1128
rect 274 1088 278 1091
rect 222 1068 230 1071
rect 222 941 225 1068
rect 310 1062 313 1148
rect 530 1138 534 1141
rect 366 1092 369 1138
rect 382 1122 385 1138
rect 250 1058 254 1061
rect 230 951 233 1058
rect 350 1052 353 1078
rect 366 1072 369 1078
rect 414 1072 417 1138
rect 462 1132 465 1138
rect 430 1082 433 1118
rect 466 1058 470 1061
rect 422 1052 425 1058
rect 414 1022 417 1048
rect 430 1032 433 1048
rect 392 1003 394 1007
rect 398 1003 401 1007
rect 405 1003 408 1007
rect 298 988 302 991
rect 262 982 265 988
rect 238 962 241 968
rect 258 958 262 961
rect 286 952 289 968
rect 294 962 297 988
rect 230 948 238 951
rect 222 938 230 941
rect 238 872 241 948
rect 390 942 393 978
rect 430 931 433 1028
rect 438 962 441 988
rect 478 982 481 1138
rect 494 1132 497 1138
rect 542 1122 545 1528
rect 630 1492 633 1538
rect 702 1492 705 1638
rect 710 1562 713 1588
rect 726 1562 729 1568
rect 742 1562 745 1648
rect 758 1642 761 1668
rect 774 1661 777 1668
rect 766 1658 777 1661
rect 782 1662 785 1728
rect 754 1618 758 1621
rect 766 1602 769 1658
rect 762 1588 766 1591
rect 770 1568 774 1571
rect 746 1558 750 1561
rect 782 1552 785 1658
rect 790 1652 793 1658
rect 798 1652 801 1688
rect 806 1672 809 1818
rect 822 1742 825 1858
rect 830 1832 833 1858
rect 830 1752 833 1818
rect 846 1752 849 1778
rect 862 1742 865 1858
rect 870 1822 873 1858
rect 894 1852 897 1858
rect 910 1832 913 1848
rect 886 1752 889 1768
rect 926 1752 929 1858
rect 934 1772 937 1988
rect 950 1962 953 1968
rect 966 1952 969 1968
rect 958 1892 961 1948
rect 974 1912 977 2048
rect 990 2032 993 2058
rect 1006 2012 1009 2058
rect 982 1962 985 1978
rect 1014 1972 1017 2058
rect 1022 1992 1025 2228
rect 1030 2132 1033 2148
rect 1038 2142 1041 2218
rect 1046 2142 1049 2208
rect 1054 2132 1057 2148
rect 1030 2062 1033 2128
rect 1038 2072 1041 2108
rect 1062 2102 1065 2218
rect 1070 2192 1073 2228
rect 1070 2152 1073 2168
rect 1086 2142 1089 2228
rect 1094 2142 1097 2248
rect 1126 2161 1129 2348
rect 1150 2342 1153 2408
rect 1182 2392 1185 2398
rect 1178 2368 1182 2371
rect 1158 2362 1161 2368
rect 1162 2348 1166 2351
rect 1138 2338 1142 2341
rect 1174 2322 1177 2368
rect 1206 2342 1209 2418
rect 1214 2352 1217 2478
rect 1238 2462 1241 2518
rect 1270 2472 1273 2488
rect 1278 2472 1281 2548
rect 1286 2482 1289 2548
rect 1326 2541 1329 2618
rect 1416 2603 1418 2607
rect 1422 2603 1425 2607
rect 1429 2603 1432 2607
rect 1342 2560 1345 2579
rect 1334 2552 1337 2558
rect 1326 2538 1337 2541
rect 1294 2492 1297 2528
rect 1334 2482 1337 2538
rect 1374 2511 1377 2538
rect 1390 2532 1393 2578
rect 1430 2542 1433 2548
rect 1374 2508 1385 2511
rect 1382 2492 1385 2508
rect 1454 2492 1457 2668
rect 1470 2622 1473 2748
rect 1478 2682 1481 2748
rect 1478 2662 1481 2668
rect 1406 2472 1409 2488
rect 1462 2482 1465 2488
rect 1370 2468 1374 2471
rect 1270 2442 1273 2468
rect 1278 2462 1281 2468
rect 1430 2462 1433 2468
rect 1438 2462 1441 2478
rect 1470 2472 1473 2618
rect 1486 2532 1489 2708
rect 1558 2702 1561 2748
rect 1614 2732 1617 2738
rect 1526 2672 1529 2678
rect 1542 2672 1545 2678
rect 1582 2662 1585 2698
rect 1494 2622 1497 2650
rect 1542 2592 1545 2648
rect 1518 2552 1521 2558
rect 1502 2532 1505 2538
rect 1486 2472 1489 2528
rect 1518 2512 1521 2518
rect 1518 2472 1521 2508
rect 1534 2492 1537 2568
rect 1354 2458 1358 2461
rect 1370 2458 1374 2461
rect 1306 2438 1310 2441
rect 1230 2412 1233 2418
rect 1222 2360 1225 2379
rect 1310 2372 1313 2438
rect 1318 2432 1321 2458
rect 1326 2452 1329 2458
rect 1346 2448 1350 2451
rect 1318 2352 1321 2428
rect 1206 2282 1209 2338
rect 1214 2302 1217 2348
rect 1254 2332 1257 2338
rect 1270 2332 1273 2338
rect 1318 2312 1321 2338
rect 1190 2262 1193 2268
rect 1246 2262 1249 2298
rect 1318 2292 1321 2308
rect 1334 2292 1337 2418
rect 1342 2362 1345 2418
rect 1350 2392 1353 2398
rect 1306 2268 1310 2271
rect 1158 2231 1161 2250
rect 1154 2188 1158 2191
rect 1122 2158 1129 2161
rect 1110 2152 1113 2158
rect 1118 2142 1121 2148
rect 1046 2062 1049 2068
rect 1054 2062 1057 2098
rect 1062 2092 1065 2098
rect 1070 2092 1073 2128
rect 1078 2112 1081 2138
rect 1142 2122 1145 2138
rect 1102 2062 1105 2068
rect 1074 2058 1078 2061
rect 1030 2032 1033 2058
rect 1030 2012 1033 2018
rect 1054 2002 1057 2058
rect 1062 2048 1070 2051
rect 1014 1962 1017 1968
rect 998 1952 1001 1958
rect 1030 1952 1033 1968
rect 982 1942 985 1948
rect 1022 1942 1025 1948
rect 1002 1938 1006 1941
rect 974 1892 977 1898
rect 1006 1872 1009 1878
rect 962 1868 966 1871
rect 986 1858 990 1861
rect 958 1812 961 1848
rect 954 1768 958 1771
rect 910 1742 913 1748
rect 866 1738 870 1741
rect 814 1702 817 1718
rect 830 1692 833 1738
rect 838 1732 841 1738
rect 918 1732 921 1748
rect 818 1658 822 1661
rect 822 1648 830 1651
rect 814 1562 817 1568
rect 762 1548 766 1551
rect 742 1532 745 1548
rect 814 1542 817 1548
rect 782 1502 785 1538
rect 566 1462 569 1478
rect 630 1472 633 1488
rect 670 1472 673 1478
rect 718 1472 721 1478
rect 798 1472 801 1478
rect 650 1468 654 1471
rect 754 1468 758 1471
rect 726 1462 729 1468
rect 602 1458 606 1461
rect 642 1458 646 1461
rect 746 1458 750 1461
rect 786 1458 790 1461
rect 550 1432 553 1448
rect 558 1442 561 1448
rect 566 1432 569 1448
rect 590 1442 593 1448
rect 574 1402 577 1438
rect 598 1432 601 1438
rect 606 1402 609 1438
rect 646 1432 649 1458
rect 574 1332 577 1338
rect 590 1292 593 1328
rect 550 1252 553 1278
rect 562 1258 566 1261
rect 570 1238 574 1241
rect 558 1212 561 1218
rect 550 1162 553 1178
rect 558 1142 561 1198
rect 574 1172 577 1238
rect 582 1232 585 1268
rect 590 1262 593 1278
rect 654 1272 657 1458
rect 678 1442 681 1448
rect 686 1432 689 1458
rect 798 1442 801 1468
rect 686 1392 689 1418
rect 686 1372 689 1388
rect 670 1342 673 1368
rect 670 1338 671 1342
rect 675 1338 678 1341
rect 662 1272 665 1288
rect 618 1268 622 1271
rect 630 1262 633 1268
rect 602 1258 606 1261
rect 614 1252 617 1258
rect 614 1192 617 1208
rect 586 1178 590 1181
rect 566 1162 569 1168
rect 574 1122 577 1158
rect 582 1152 585 1168
rect 630 1152 633 1248
rect 638 1222 641 1268
rect 670 1262 673 1268
rect 678 1262 681 1328
rect 686 1282 689 1298
rect 694 1292 697 1438
rect 806 1422 809 1518
rect 822 1492 825 1648
rect 838 1642 841 1668
rect 846 1662 849 1698
rect 862 1692 865 1718
rect 870 1682 873 1718
rect 918 1712 921 1718
rect 896 1703 898 1707
rect 902 1703 905 1707
rect 909 1703 912 1707
rect 882 1658 886 1661
rect 894 1652 897 1678
rect 926 1662 929 1748
rect 934 1722 937 1748
rect 942 1742 945 1748
rect 950 1732 953 1738
rect 966 1692 969 1858
rect 974 1832 977 1858
rect 998 1841 1001 1868
rect 1014 1862 1017 1888
rect 1038 1882 1041 1998
rect 1062 1992 1065 2048
rect 1110 2042 1113 2048
rect 1054 1952 1057 1968
rect 1070 1962 1073 1968
rect 1070 1952 1073 1958
rect 1062 1892 1065 1948
rect 1078 1942 1081 1988
rect 1086 1952 1089 2028
rect 1102 1952 1105 1978
rect 1090 1948 1097 1951
rect 1086 1932 1089 1938
rect 1038 1872 1041 1878
rect 1094 1872 1097 1948
rect 1118 1941 1121 2108
rect 1134 2072 1137 2088
rect 1126 2052 1129 2058
rect 1142 2042 1145 2048
rect 1126 2032 1129 2038
rect 1150 2022 1153 2058
rect 1158 2042 1161 2048
rect 1158 2012 1161 2038
rect 1114 1938 1121 1941
rect 1042 1858 1046 1861
rect 1074 1858 1078 1861
rect 990 1838 1001 1841
rect 990 1742 993 1838
rect 1030 1832 1033 1848
rect 998 1792 1001 1828
rect 978 1688 982 1691
rect 942 1672 945 1688
rect 954 1668 961 1671
rect 906 1658 910 1661
rect 930 1658 934 1661
rect 918 1652 921 1658
rect 950 1652 953 1658
rect 878 1632 881 1638
rect 830 1552 833 1618
rect 814 1462 817 1468
rect 822 1432 825 1438
rect 830 1431 833 1548
rect 838 1542 841 1578
rect 846 1562 849 1588
rect 886 1582 889 1598
rect 866 1548 870 1551
rect 846 1502 849 1518
rect 854 1492 857 1498
rect 838 1472 841 1478
rect 862 1472 865 1548
rect 878 1542 881 1578
rect 886 1552 889 1578
rect 894 1562 897 1648
rect 958 1642 961 1668
rect 982 1662 985 1668
rect 974 1642 977 1648
rect 906 1588 910 1591
rect 942 1572 945 1638
rect 942 1552 945 1568
rect 958 1552 961 1578
rect 898 1548 902 1551
rect 962 1548 966 1551
rect 974 1542 977 1548
rect 870 1532 873 1538
rect 870 1512 873 1518
rect 870 1462 873 1508
rect 896 1503 898 1507
rect 902 1503 905 1507
rect 909 1503 912 1507
rect 878 1472 881 1478
rect 906 1468 910 1471
rect 878 1452 881 1458
rect 846 1432 849 1448
rect 886 1442 889 1468
rect 918 1442 921 1538
rect 926 1472 929 1488
rect 830 1428 841 1431
rect 726 1351 729 1418
rect 758 1391 761 1408
rect 766 1402 769 1418
rect 758 1388 766 1391
rect 750 1362 753 1378
rect 782 1362 785 1408
rect 798 1372 801 1378
rect 806 1372 809 1398
rect 718 1348 729 1351
rect 830 1361 833 1418
rect 826 1358 833 1361
rect 734 1352 737 1358
rect 790 1352 793 1358
rect 838 1352 841 1428
rect 862 1392 865 1408
rect 846 1362 849 1378
rect 858 1368 862 1371
rect 802 1348 806 1351
rect 826 1348 830 1351
rect 702 1342 705 1348
rect 710 1342 713 1348
rect 702 1282 705 1338
rect 718 1302 721 1348
rect 754 1338 758 1341
rect 710 1262 713 1268
rect 650 1248 654 1251
rect 662 1242 665 1248
rect 710 1242 713 1248
rect 646 1172 649 1178
rect 606 1132 609 1138
rect 518 1082 521 1118
rect 550 1102 553 1118
rect 534 1082 537 1088
rect 518 1052 521 1068
rect 486 1031 489 1050
rect 534 1012 537 1078
rect 606 1072 609 1128
rect 614 1092 617 1108
rect 482 968 486 971
rect 614 960 617 979
rect 438 942 441 948
rect 526 942 529 948
rect 582 942 585 948
rect 622 942 625 948
rect 430 928 441 931
rect 374 922 377 928
rect 438 882 441 928
rect 262 872 265 878
rect 222 868 230 871
rect 214 692 217 728
rect 222 712 225 868
rect 238 862 241 868
rect 254 852 257 858
rect 238 842 241 848
rect 230 742 233 778
rect 302 751 305 868
rect 314 768 318 771
rect 326 762 329 838
rect 302 748 310 751
rect 290 738 294 741
rect 230 692 233 738
rect 270 672 273 738
rect 302 712 305 738
rect 310 702 313 748
rect 334 742 337 868
rect 362 838 366 841
rect 392 803 394 807
rect 398 803 401 807
rect 405 803 408 807
rect 390 782 393 788
rect 426 778 430 781
rect 338 738 342 741
rect 366 682 369 738
rect 438 712 441 878
rect 454 872 457 878
rect 510 862 513 938
rect 566 902 569 928
rect 554 868 558 871
rect 454 702 457 858
rect 550 852 553 858
rect 558 852 561 868
rect 486 831 489 850
rect 534 812 537 818
rect 470 702 473 748
rect 526 742 529 748
rect 566 742 569 898
rect 618 888 622 891
rect 630 871 633 1148
rect 638 1142 641 1158
rect 646 1132 649 1148
rect 654 1082 657 1218
rect 694 1202 697 1238
rect 726 1212 729 1338
rect 742 1332 745 1338
rect 742 1272 745 1318
rect 750 1292 753 1308
rect 758 1282 761 1318
rect 766 1312 769 1348
rect 790 1302 793 1348
rect 846 1342 849 1358
rect 822 1292 825 1308
rect 838 1292 841 1328
rect 854 1302 857 1358
rect 862 1352 865 1358
rect 770 1288 774 1291
rect 734 1262 737 1268
rect 698 1158 702 1161
rect 662 1082 665 1158
rect 682 1148 686 1151
rect 714 1148 718 1151
rect 702 1142 705 1148
rect 670 1132 673 1138
rect 670 1102 673 1128
rect 642 1068 646 1071
rect 638 942 641 1068
rect 654 1062 657 1068
rect 646 892 649 1058
rect 678 1052 681 1118
rect 686 1062 689 1138
rect 714 1118 718 1121
rect 726 1072 729 1148
rect 734 1112 737 1238
rect 742 1142 745 1228
rect 750 1172 753 1218
rect 766 1152 769 1198
rect 750 1132 753 1148
rect 774 1142 777 1168
rect 766 1072 769 1118
rect 738 1068 742 1071
rect 746 1058 750 1061
rect 718 1052 721 1058
rect 658 1048 662 1051
rect 706 1048 710 1051
rect 770 1048 774 1051
rect 662 992 665 1038
rect 670 1022 673 1048
rect 666 938 670 941
rect 654 932 657 938
rect 622 868 633 871
rect 574 762 577 788
rect 382 672 385 678
rect 186 658 190 661
rect 182 622 185 648
rect 198 592 201 668
rect 326 662 329 668
rect 150 552 153 558
rect 186 548 190 551
rect 174 542 177 548
rect 142 532 145 538
rect 182 462 185 468
rect 166 422 169 450
rect 110 262 113 268
rect 58 188 62 191
rect 78 142 81 188
rect 142 142 145 318
rect 150 262 153 348
rect 190 332 193 528
rect 214 392 217 618
rect 230 552 233 658
rect 414 622 417 650
rect 282 618 286 621
rect 392 603 394 607
rect 398 603 401 607
rect 405 603 408 607
rect 246 560 249 579
rect 230 462 233 548
rect 278 542 281 578
rect 406 562 409 568
rect 422 552 425 698
rect 438 662 441 698
rect 470 672 473 678
rect 438 552 441 558
rect 426 548 430 551
rect 470 542 473 668
rect 426 538 430 541
rect 294 522 297 528
rect 286 482 289 488
rect 398 472 401 528
rect 270 462 273 468
rect 222 422 225 448
rect 254 362 257 388
rect 302 352 305 358
rect 326 352 329 458
rect 406 442 409 518
rect 370 428 374 431
rect 392 403 394 407
rect 398 403 401 407
rect 405 403 408 407
rect 358 360 361 379
rect 258 348 262 351
rect 338 348 342 351
rect 278 342 281 348
rect 390 342 393 368
rect 206 332 209 338
rect 190 302 193 328
rect 262 282 265 288
rect 194 258 198 261
rect 158 222 161 248
rect 166 152 169 258
rect 214 222 217 250
rect 246 242 249 268
rect 358 252 361 308
rect 406 302 409 328
rect 374 262 377 288
rect 454 272 457 518
rect 470 472 473 538
rect 478 392 481 708
rect 510 672 513 728
rect 534 672 537 688
rect 542 552 545 558
rect 550 541 553 618
rect 558 592 561 728
rect 582 552 585 808
rect 614 792 617 808
rect 598 752 601 758
rect 622 752 625 868
rect 654 862 657 928
rect 662 872 665 938
rect 678 912 681 1048
rect 750 1042 753 1048
rect 698 1038 702 1041
rect 714 1018 718 1021
rect 686 961 689 1018
rect 726 982 729 1038
rect 782 992 785 1258
rect 790 1192 793 1268
rect 830 1262 833 1268
rect 798 1192 801 1258
rect 822 1252 825 1258
rect 838 1252 841 1258
rect 790 1162 793 1188
rect 798 1082 801 1188
rect 814 1181 817 1218
rect 814 1178 825 1181
rect 806 1142 809 1148
rect 814 1142 817 1168
rect 822 1152 825 1178
rect 838 1162 841 1238
rect 846 1142 849 1248
rect 854 1212 857 1268
rect 862 1262 865 1338
rect 870 1272 873 1428
rect 894 1412 897 1418
rect 898 1358 902 1361
rect 914 1358 918 1361
rect 922 1348 926 1351
rect 934 1351 937 1468
rect 942 1362 945 1368
rect 934 1348 945 1351
rect 894 1342 897 1348
rect 886 1292 889 1338
rect 934 1322 937 1338
rect 896 1303 898 1307
rect 902 1303 905 1307
rect 909 1303 912 1307
rect 942 1292 945 1348
rect 886 1272 889 1278
rect 942 1272 945 1288
rect 950 1281 953 1538
rect 966 1532 969 1538
rect 958 1362 961 1508
rect 982 1492 985 1568
rect 990 1512 993 1728
rect 1006 1671 1009 1758
rect 1014 1722 1017 1818
rect 1022 1752 1025 1758
rect 1054 1752 1057 1858
rect 1062 1822 1065 1848
rect 1022 1731 1025 1748
rect 1046 1742 1049 1748
rect 1034 1738 1038 1741
rect 1054 1732 1057 1738
rect 1022 1728 1033 1731
rect 1006 1668 1014 1671
rect 1002 1658 1006 1661
rect 1006 1632 1009 1658
rect 974 1442 977 1468
rect 986 1458 990 1461
rect 986 1448 990 1451
rect 966 1342 969 1438
rect 966 1292 969 1308
rect 974 1302 977 1318
rect 950 1278 961 1281
rect 930 1268 934 1271
rect 870 1172 873 1268
rect 878 1262 881 1268
rect 910 1232 913 1268
rect 950 1262 953 1268
rect 938 1258 945 1261
rect 918 1222 921 1258
rect 942 1192 945 1258
rect 918 1172 921 1178
rect 926 1172 929 1178
rect 858 1158 862 1161
rect 942 1158 950 1161
rect 958 1161 961 1278
rect 982 1272 985 1418
rect 998 1282 1001 1598
rect 1006 1542 1009 1548
rect 1014 1542 1017 1668
rect 1022 1652 1025 1658
rect 1022 1602 1025 1648
rect 1030 1562 1033 1728
rect 1038 1692 1041 1718
rect 1062 1692 1065 1768
rect 1078 1762 1081 1818
rect 1078 1732 1081 1758
rect 1094 1752 1097 1858
rect 1102 1851 1105 1908
rect 1110 1882 1113 1938
rect 1118 1912 1121 1928
rect 1114 1858 1118 1861
rect 1102 1848 1113 1851
rect 1102 1822 1105 1828
rect 1110 1792 1113 1848
rect 1126 1842 1129 2008
rect 1158 1972 1161 2008
rect 1174 1992 1177 2208
rect 1246 2152 1249 2258
rect 1318 2252 1321 2278
rect 1342 2262 1345 2348
rect 1358 2342 1361 2358
rect 1318 2232 1321 2248
rect 1282 2218 1286 2221
rect 1182 2072 1185 2078
rect 1190 2062 1193 2148
rect 1230 2132 1233 2138
rect 1246 2132 1249 2138
rect 1230 2102 1233 2128
rect 1198 2072 1201 2098
rect 1206 2061 1209 2088
rect 1286 2082 1289 2198
rect 1294 2162 1297 2188
rect 1318 2152 1321 2158
rect 1314 2138 1318 2141
rect 1270 2072 1273 2078
rect 1202 2058 1209 2061
rect 1218 2058 1222 2061
rect 1162 1958 1166 1961
rect 1134 1952 1137 1958
rect 1170 1948 1174 1951
rect 1146 1938 1150 1941
rect 1162 1938 1166 1941
rect 1158 1872 1161 1888
rect 1170 1868 1174 1871
rect 1146 1858 1150 1861
rect 1182 1861 1185 1978
rect 1190 1892 1193 2048
rect 1238 2031 1241 2050
rect 1230 1962 1233 2018
rect 1262 1982 1265 1988
rect 1250 1968 1254 1971
rect 1262 1962 1265 1968
rect 1234 1958 1249 1961
rect 1210 1948 1214 1951
rect 1238 1942 1241 1948
rect 1198 1932 1201 1938
rect 1198 1872 1201 1928
rect 1222 1912 1225 1918
rect 1238 1882 1241 1918
rect 1214 1872 1217 1878
rect 1178 1858 1185 1861
rect 1210 1858 1222 1861
rect 1134 1842 1137 1848
rect 1126 1772 1129 1838
rect 1134 1822 1137 1838
rect 1150 1792 1153 1858
rect 1106 1768 1110 1771
rect 1138 1758 1142 1761
rect 1150 1752 1153 1758
rect 1070 1692 1073 1718
rect 1094 1682 1097 1748
rect 1118 1742 1121 1748
rect 1102 1682 1105 1708
rect 1142 1672 1145 1708
rect 1166 1692 1169 1828
rect 1182 1792 1185 1858
rect 1246 1852 1249 1958
rect 1254 1862 1257 1878
rect 1194 1848 1201 1851
rect 1198 1792 1201 1848
rect 1222 1842 1225 1848
rect 1222 1792 1225 1808
rect 1226 1788 1230 1791
rect 1230 1772 1233 1778
rect 1186 1768 1190 1771
rect 1246 1762 1249 1848
rect 1262 1842 1265 1958
rect 1270 1942 1273 2058
rect 1302 1972 1305 1978
rect 1278 1952 1281 1958
rect 1310 1951 1313 1968
rect 1318 1962 1321 1978
rect 1306 1948 1313 1951
rect 1326 1952 1329 2238
rect 1334 2132 1337 2138
rect 1342 2082 1345 2248
rect 1366 2242 1369 2438
rect 1374 2352 1377 2448
rect 1382 2422 1385 2448
rect 1398 2392 1401 2458
rect 1454 2422 1457 2448
rect 1416 2403 1418 2407
rect 1422 2403 1425 2407
rect 1429 2403 1432 2407
rect 1438 2372 1441 2408
rect 1454 2362 1457 2368
rect 1386 2348 1390 2351
rect 1462 2342 1465 2398
rect 1470 2352 1473 2458
rect 1502 2452 1505 2458
rect 1490 2448 1494 2451
rect 1502 2441 1505 2448
rect 1494 2438 1505 2441
rect 1514 2438 1518 2441
rect 1494 2432 1497 2438
rect 1502 2422 1505 2428
rect 1478 2392 1481 2418
rect 1526 2412 1529 2468
rect 1542 2452 1545 2548
rect 1558 2522 1561 2558
rect 1574 2542 1577 2548
rect 1582 2542 1585 2608
rect 1598 2532 1601 2728
rect 1686 2692 1689 2748
rect 1626 2688 1630 2691
rect 1646 2672 1649 2678
rect 1658 2668 1662 2671
rect 1694 2662 1697 2748
rect 1742 2701 1745 2808
rect 1774 2802 1777 2848
rect 1782 2832 1785 2858
rect 1790 2842 1793 2858
rect 1754 2748 1758 2751
rect 1814 2732 1817 2738
rect 1798 2722 1801 2728
rect 1742 2698 1753 2701
rect 1750 2682 1753 2698
rect 1734 2672 1737 2678
rect 1634 2648 1638 2651
rect 1654 2612 1657 2658
rect 1702 2631 1705 2650
rect 1622 2560 1625 2579
rect 1750 2572 1753 2678
rect 1846 2672 1849 2848
rect 1858 2828 1862 2831
rect 1862 2762 1865 2788
rect 1870 2752 1873 2778
rect 1878 2662 1881 2808
rect 1886 2782 1889 2858
rect 1902 2831 1905 2850
rect 1998 2822 2001 3128
rect 2022 3092 2025 3128
rect 2046 3092 2049 3128
rect 2058 3058 2065 3061
rect 2030 2992 2033 3058
rect 2062 3042 2065 3058
rect 2038 2922 2041 2938
rect 2038 2912 2041 2918
rect 2030 2892 2033 2898
rect 2046 2882 2049 2988
rect 2054 2902 2057 2948
rect 2062 2942 2065 3038
rect 2070 2992 2073 3128
rect 2142 3128 2146 3132
rect 2174 3128 2178 3132
rect 2246 3128 2250 3132
rect 2406 3128 2410 3132
rect 2486 3128 2490 3132
rect 2566 3128 2570 3132
rect 2638 3128 2642 3132
rect 2142 3102 2145 3128
rect 2174 3102 2177 3128
rect 2086 3062 2089 3068
rect 2130 3058 2134 3061
rect 2090 3018 2094 3021
rect 2082 2988 2086 2991
rect 2126 2952 2129 3058
rect 2174 3012 2177 3078
rect 2190 2992 2193 3068
rect 2222 3031 2225 3050
rect 2230 2962 2233 2988
rect 2086 2892 2089 2948
rect 2182 2942 2185 2948
rect 2166 2922 2169 2928
rect 2174 2882 2177 2908
rect 2158 2862 2161 2868
rect 2214 2862 2217 2948
rect 2070 2832 2073 2858
rect 2074 2828 2081 2831
rect 1886 2662 1889 2768
rect 2054 2762 2057 2788
rect 2078 2762 2081 2828
rect 2086 2792 2089 2848
rect 2094 2762 2097 2768
rect 1990 2732 1993 2758
rect 2090 2748 2094 2751
rect 2006 2732 2009 2738
rect 2054 2732 2057 2748
rect 2102 2732 2105 2858
rect 2126 2822 2129 2850
rect 2214 2772 2217 2858
rect 2210 2758 2217 2761
rect 2134 2752 2137 2758
rect 2162 2748 2166 2751
rect 1910 2672 1913 2718
rect 1928 2703 1930 2707
rect 1934 2703 1937 2707
rect 1941 2703 1944 2707
rect 1926 2682 1929 2688
rect 2046 2672 2049 2678
rect 1906 2658 1910 2661
rect 1854 2642 1857 2648
rect 1766 2592 1769 2608
rect 1610 2548 1614 2551
rect 1755 2548 1758 2551
rect 1774 2542 1777 2548
rect 1782 2542 1785 2578
rect 1806 2572 1809 2618
rect 1822 2572 1825 2608
rect 1830 2552 1833 2558
rect 1838 2552 1841 2638
rect 1850 2588 1854 2591
rect 1878 2552 1881 2658
rect 1886 2552 1889 2658
rect 1894 2582 1897 2618
rect 1894 2552 1897 2558
rect 1942 2552 1945 2558
rect 1822 2548 1830 2551
rect 1654 2512 1657 2538
rect 1670 2522 1673 2528
rect 1630 2492 1633 2508
rect 1666 2488 1670 2491
rect 1734 2482 1737 2488
rect 1766 2482 1769 2528
rect 1790 2502 1793 2518
rect 1722 2478 1726 2481
rect 1678 2472 1681 2478
rect 1626 2468 1630 2471
rect 1582 2452 1585 2458
rect 1598 2452 1601 2468
rect 1646 2462 1649 2468
rect 1654 2462 1657 2468
rect 1614 2452 1617 2458
rect 1630 2442 1633 2448
rect 1646 2442 1649 2458
rect 1570 2438 1574 2441
rect 1550 2432 1553 2438
rect 1582 2432 1585 2438
rect 1662 2432 1665 2448
rect 1526 2352 1529 2388
rect 1490 2348 1494 2351
rect 1538 2348 1542 2351
rect 1386 2338 1390 2341
rect 1402 2338 1406 2341
rect 1546 2338 1550 2341
rect 1382 2212 1385 2338
rect 1390 2262 1393 2298
rect 1390 2222 1393 2248
rect 1350 2022 1353 2158
rect 1358 2132 1361 2148
rect 1366 2142 1369 2168
rect 1382 2162 1385 2168
rect 1366 2101 1369 2138
rect 1390 2132 1393 2188
rect 1398 2182 1401 2338
rect 1398 2152 1401 2178
rect 1406 2112 1409 2318
rect 1438 2282 1441 2338
rect 1478 2332 1481 2338
rect 1446 2302 1449 2318
rect 1454 2282 1457 2318
rect 1494 2312 1497 2338
rect 1502 2332 1505 2338
rect 1510 2292 1513 2318
rect 1416 2203 1418 2207
rect 1422 2203 1425 2207
rect 1429 2203 1432 2207
rect 1426 2158 1430 2161
rect 1414 2132 1417 2138
rect 1438 2112 1441 2268
rect 1518 2262 1521 2338
rect 1366 2098 1377 2101
rect 1362 2048 1366 2051
rect 1342 1972 1345 1978
rect 1374 1962 1377 2098
rect 1446 2092 1449 2218
rect 1494 2202 1497 2258
rect 1518 2222 1521 2258
rect 1542 2222 1545 2328
rect 1582 2292 1585 2418
rect 1638 2392 1641 2428
rect 1686 2412 1689 2468
rect 1694 2462 1697 2478
rect 1702 2472 1705 2478
rect 1798 2472 1801 2498
rect 1806 2492 1809 2538
rect 1814 2512 1817 2518
rect 1714 2468 1718 2471
rect 1710 2432 1713 2458
rect 1742 2442 1745 2468
rect 1750 2462 1753 2468
rect 1806 2452 1809 2488
rect 1822 2462 1825 2548
rect 1870 2522 1873 2528
rect 1870 2482 1873 2488
rect 1830 2462 1833 2468
rect 1858 2458 1862 2461
rect 1774 2442 1777 2448
rect 1646 2368 1654 2371
rect 1646 2352 1649 2368
rect 1654 2352 1657 2358
rect 1666 2348 1670 2351
rect 1678 2342 1681 2398
rect 1742 2392 1745 2428
rect 1690 2358 1694 2361
rect 1710 2352 1713 2358
rect 1722 2348 1726 2351
rect 1734 2342 1737 2388
rect 1750 2372 1753 2408
rect 1758 2402 1761 2418
rect 1774 2372 1777 2438
rect 1782 2362 1785 2418
rect 1798 2392 1801 2428
rect 1806 2382 1809 2418
rect 1790 2362 1793 2368
rect 1806 2362 1809 2368
rect 1750 2352 1753 2358
rect 1778 2348 1782 2351
rect 1650 2338 1654 2341
rect 1698 2338 1702 2341
rect 1606 2322 1609 2328
rect 1622 2322 1625 2328
rect 1622 2288 1638 2291
rect 1550 2252 1553 2278
rect 1590 2272 1593 2278
rect 1598 2262 1601 2288
rect 1622 2282 1625 2288
rect 1610 2278 1614 2281
rect 1606 2262 1609 2268
rect 1566 2242 1569 2258
rect 1606 2232 1609 2258
rect 1630 2252 1633 2268
rect 1638 2262 1641 2278
rect 1534 2212 1537 2218
rect 1462 2162 1465 2188
rect 1510 2152 1513 2198
rect 1486 2092 1489 2108
rect 1382 2072 1385 2078
rect 1406 2072 1409 2078
rect 1494 2072 1497 2098
rect 1462 2062 1465 2068
rect 1470 2062 1473 2068
rect 1382 2042 1385 2048
rect 1398 2032 1401 2058
rect 1406 2011 1409 2058
rect 1398 2008 1409 2011
rect 1390 1992 1393 1998
rect 1382 1952 1385 1988
rect 1362 1948 1369 1951
rect 1326 1942 1329 1948
rect 1354 1938 1358 1941
rect 1278 1932 1281 1938
rect 1354 1928 1358 1931
rect 1310 1892 1313 1908
rect 1334 1882 1337 1918
rect 1294 1872 1297 1878
rect 1342 1872 1345 1928
rect 1366 1892 1369 1948
rect 1270 1868 1278 1871
rect 1330 1868 1334 1871
rect 1270 1862 1273 1868
rect 1282 1858 1286 1861
rect 1354 1858 1358 1861
rect 1302 1852 1305 1858
rect 1314 1848 1321 1851
rect 1254 1832 1257 1838
rect 1262 1832 1265 1838
rect 1318 1792 1321 1848
rect 1282 1788 1297 1791
rect 1262 1762 1265 1788
rect 1198 1752 1201 1758
rect 1174 1742 1177 1748
rect 1198 1742 1201 1748
rect 1206 1732 1209 1758
rect 1270 1752 1273 1788
rect 1274 1748 1278 1751
rect 1286 1742 1289 1778
rect 1294 1762 1297 1788
rect 1326 1782 1329 1858
rect 1366 1842 1369 1848
rect 1306 1768 1310 1771
rect 1302 1752 1305 1758
rect 1334 1752 1337 1828
rect 1350 1822 1353 1828
rect 1346 1748 1350 1751
rect 1250 1738 1254 1741
rect 1178 1678 1182 1681
rect 1042 1668 1046 1671
rect 1202 1668 1206 1671
rect 1046 1662 1049 1668
rect 1086 1652 1089 1658
rect 1038 1642 1041 1648
rect 1070 1642 1073 1648
rect 1094 1642 1097 1668
rect 1214 1662 1217 1738
rect 1230 1692 1233 1728
rect 1246 1672 1249 1718
rect 1262 1692 1265 1728
rect 1294 1692 1297 1748
rect 1358 1742 1361 1828
rect 1374 1822 1377 1868
rect 1382 1832 1385 1938
rect 1390 1932 1393 1938
rect 1390 1852 1393 1908
rect 1390 1832 1393 1848
rect 1390 1821 1393 1828
rect 1382 1818 1393 1821
rect 1374 1802 1377 1818
rect 1382 1752 1385 1818
rect 1398 1752 1401 2008
rect 1416 2003 1418 2007
rect 1422 2003 1425 2007
rect 1429 2003 1432 2007
rect 1438 1991 1441 2028
rect 1430 1988 1441 1991
rect 1430 1952 1433 1988
rect 1438 1952 1441 1958
rect 1462 1942 1465 2008
rect 1486 1992 1489 2048
rect 1470 1952 1473 1978
rect 1442 1938 1446 1941
rect 1406 1912 1409 1938
rect 1462 1932 1465 1938
rect 1446 1892 1449 1908
rect 1454 1882 1457 1918
rect 1478 1912 1481 1958
rect 1486 1932 1489 1948
rect 1494 1911 1497 1968
rect 1486 1908 1497 1911
rect 1478 1892 1481 1898
rect 1406 1862 1409 1878
rect 1470 1872 1473 1878
rect 1462 1852 1465 1858
rect 1470 1848 1478 1851
rect 1446 1842 1449 1848
rect 1418 1838 1422 1841
rect 1406 1812 1409 1818
rect 1416 1803 1418 1807
rect 1422 1803 1425 1807
rect 1429 1803 1432 1807
rect 1438 1772 1441 1808
rect 1470 1792 1473 1848
rect 1486 1812 1489 1908
rect 1502 1872 1505 2058
rect 1510 1902 1513 2138
rect 1526 2132 1529 2138
rect 1526 1952 1529 2078
rect 1534 1892 1537 2098
rect 1566 2082 1569 2148
rect 1598 2082 1601 2088
rect 1606 2072 1609 2208
rect 1646 2192 1649 2328
rect 1662 2272 1665 2278
rect 1670 2272 1673 2338
rect 1694 2312 1697 2328
rect 1670 2262 1673 2268
rect 1678 2262 1681 2298
rect 1710 2292 1713 2298
rect 1718 2282 1721 2338
rect 1758 2332 1761 2348
rect 1766 2332 1769 2338
rect 1726 2282 1729 2318
rect 1750 2302 1753 2328
rect 1702 2272 1705 2278
rect 1774 2272 1777 2308
rect 1730 2268 1734 2271
rect 1754 2258 1758 2261
rect 1618 2148 1622 2151
rect 1630 2142 1633 2188
rect 1654 2152 1657 2198
rect 1662 2192 1665 2258
rect 1694 2252 1697 2258
rect 1782 2252 1785 2258
rect 1682 2238 1686 2241
rect 1758 2232 1761 2248
rect 1686 2162 1689 2168
rect 1694 2152 1697 2208
rect 1742 2152 1745 2168
rect 1766 2162 1769 2218
rect 1782 2172 1785 2228
rect 1798 2162 1801 2348
rect 1806 2282 1809 2358
rect 1814 2352 1817 2358
rect 1822 2342 1825 2428
rect 1830 2392 1833 2398
rect 1814 2282 1817 2328
rect 1814 2242 1817 2268
rect 1830 2232 1833 2358
rect 1838 2332 1841 2418
rect 1878 2352 1881 2478
rect 1886 2472 1889 2548
rect 1894 2462 1897 2548
rect 1914 2538 1918 2541
rect 1950 2522 1953 2638
rect 1990 2532 1993 2598
rect 2006 2542 2009 2548
rect 2022 2532 2025 2538
rect 1928 2503 1930 2507
rect 1934 2503 1937 2507
rect 1941 2503 1944 2507
rect 1918 2462 1921 2498
rect 1938 2468 1942 2471
rect 1950 2462 1953 2518
rect 1958 2502 1961 2518
rect 1974 2472 1977 2528
rect 1990 2482 1993 2528
rect 2030 2522 2033 2548
rect 2038 2532 2041 2548
rect 2046 2542 2049 2658
rect 2062 2552 2065 2668
rect 2102 2662 2105 2728
rect 2110 2692 2113 2748
rect 2118 2742 2121 2748
rect 2142 2732 2145 2748
rect 2134 2662 2137 2668
rect 2142 2662 2145 2668
rect 2150 2662 2153 2748
rect 2198 2742 2201 2758
rect 2158 2728 2166 2731
rect 2158 2692 2161 2728
rect 2214 2692 2217 2758
rect 2226 2748 2230 2751
rect 2226 2738 2230 2741
rect 2230 2712 2233 2738
rect 2246 2671 2249 3128
rect 2406 3102 2409 3128
rect 2486 3102 2489 3128
rect 2510 3082 2513 3088
rect 2330 3068 2334 3071
rect 2402 3068 2406 3071
rect 2434 3018 2438 3021
rect 2270 2972 2273 3018
rect 2274 2958 2278 2961
rect 2254 2942 2257 2958
rect 2294 2952 2297 2958
rect 2254 2792 2257 2818
rect 2262 2781 2265 2858
rect 2278 2851 2281 2918
rect 2286 2862 2289 2878
rect 2274 2848 2281 2851
rect 2294 2852 2297 2948
rect 2302 2932 2305 2938
rect 2310 2872 2313 2878
rect 2318 2872 2321 3018
rect 2342 2952 2345 3018
rect 2440 3003 2442 3007
rect 2446 3003 2449 3007
rect 2453 3003 2456 3007
rect 2470 2981 2473 3058
rect 2470 2978 2481 2981
rect 2478 2952 2481 2978
rect 2326 2902 2329 2948
rect 2398 2942 2401 2948
rect 2470 2942 2473 2948
rect 2334 2872 2337 2878
rect 2342 2831 2345 2918
rect 2414 2912 2417 2918
rect 2422 2882 2425 2898
rect 2342 2828 2350 2831
rect 2382 2822 2385 2858
rect 2438 2822 2441 2868
rect 2478 2862 2481 2948
rect 2470 2831 2473 2850
rect 2342 2802 2345 2818
rect 2254 2778 2265 2781
rect 2254 2682 2257 2778
rect 2262 2752 2265 2768
rect 2270 2760 2273 2779
rect 2302 2742 2305 2758
rect 2358 2752 2361 2818
rect 2440 2803 2442 2807
rect 2446 2803 2449 2807
rect 2453 2803 2456 2807
rect 2318 2732 2321 2738
rect 2258 2678 2262 2681
rect 2270 2672 2273 2718
rect 2358 2702 2361 2748
rect 2414 2742 2417 2798
rect 2462 2792 2465 2808
rect 2398 2712 2401 2718
rect 2318 2672 2321 2688
rect 2398 2682 2401 2688
rect 2386 2678 2390 2681
rect 2366 2672 2369 2678
rect 2406 2672 2409 2708
rect 2422 2682 2425 2718
rect 2246 2668 2254 2671
rect 2354 2668 2358 2671
rect 2430 2671 2433 2718
rect 2422 2668 2433 2671
rect 2166 2662 2169 2668
rect 2230 2662 2233 2668
rect 2302 2662 2305 2668
rect 2314 2658 2318 2661
rect 2330 2658 2334 2661
rect 2346 2658 2350 2661
rect 2094 2622 2097 2650
rect 2158 2642 2161 2648
rect 2142 2592 2145 2638
rect 2174 2622 2177 2658
rect 2190 2642 2193 2658
rect 2074 2558 2078 2561
rect 2090 2558 2094 2561
rect 2106 2558 2110 2561
rect 2158 2552 2161 2558
rect 2166 2552 2169 2598
rect 2082 2548 2086 2551
rect 2138 2548 2142 2551
rect 2054 2542 2057 2548
rect 2074 2538 2078 2541
rect 2006 2472 2009 2478
rect 2014 2462 2017 2498
rect 2038 2482 2041 2488
rect 1962 2458 1966 2461
rect 1978 2458 1982 2461
rect 2002 2458 2006 2461
rect 2022 2452 2025 2458
rect 1970 2448 1974 2451
rect 1910 2402 1913 2418
rect 1982 2392 1985 2448
rect 2030 2422 2033 2478
rect 2058 2468 2062 2471
rect 2070 2462 2073 2528
rect 2078 2512 2081 2538
rect 2106 2528 2110 2531
rect 2078 2478 2105 2481
rect 2078 2472 2081 2478
rect 2102 2472 2105 2478
rect 2050 2458 2054 2461
rect 2086 2452 2089 2458
rect 2038 2442 2041 2448
rect 2070 2442 2073 2448
rect 1990 2372 1993 2418
rect 1850 2348 1854 2351
rect 1886 2342 1889 2348
rect 1910 2342 1913 2368
rect 2006 2362 2009 2408
rect 2014 2392 2017 2408
rect 1950 2352 1953 2358
rect 1974 2352 1977 2358
rect 1938 2348 1942 2351
rect 2034 2348 2038 2351
rect 1998 2342 2001 2348
rect 2014 2338 2022 2341
rect 1854 2282 1857 2338
rect 1870 2332 1873 2338
rect 1862 2311 1865 2318
rect 1862 2308 1870 2311
rect 1878 2282 1881 2298
rect 1902 2282 1905 2318
rect 1910 2302 1913 2338
rect 1966 2332 1969 2338
rect 1928 2303 1930 2307
rect 1934 2303 1937 2307
rect 1941 2303 1944 2307
rect 1838 2262 1841 2278
rect 1862 2262 1865 2278
rect 1966 2272 1969 2308
rect 1990 2282 1993 2298
rect 1806 2162 1809 2178
rect 1814 2172 1817 2228
rect 1830 2162 1833 2218
rect 1758 2152 1761 2158
rect 1666 2148 1670 2151
rect 1802 2148 1806 2151
rect 1702 2142 1705 2148
rect 1718 2142 1721 2148
rect 1774 2142 1777 2148
rect 1846 2142 1849 2218
rect 1854 2152 1857 2258
rect 1870 2242 1873 2248
rect 1886 2212 1889 2268
rect 1898 2258 1902 2261
rect 1918 2252 1921 2268
rect 1974 2262 1977 2278
rect 2014 2272 2017 2338
rect 2022 2292 2025 2308
rect 2030 2302 2033 2338
rect 2038 2282 2041 2308
rect 1926 2252 1929 2258
rect 1942 2252 1945 2258
rect 1966 2251 1969 2258
rect 1990 2252 1993 2268
rect 2002 2258 2006 2261
rect 2026 2258 2030 2261
rect 2038 2252 2041 2268
rect 1966 2248 1977 2251
rect 2018 2248 2022 2251
rect 1910 2232 1913 2248
rect 1974 2242 1977 2248
rect 1954 2238 1958 2241
rect 1918 2162 1921 2238
rect 2046 2232 2049 2318
rect 2054 2262 2057 2368
rect 2070 2362 2073 2438
rect 2078 2351 2081 2378
rect 2074 2348 2081 2351
rect 2074 2338 2078 2341
rect 2062 2332 2065 2338
rect 1974 2162 1977 2228
rect 2006 2168 2025 2171
rect 1978 2158 1982 2161
rect 2006 2161 2009 2168
rect 1990 2158 2009 2161
rect 1966 2152 1969 2158
rect 1906 2148 1910 2151
rect 1990 2151 1993 2158
rect 1986 2148 1993 2151
rect 2002 2148 2006 2151
rect 1682 2138 1686 2141
rect 1614 2122 1617 2128
rect 1618 2068 1622 2071
rect 1590 2062 1593 2068
rect 1570 2058 1574 2061
rect 1566 2052 1569 2058
rect 1550 2002 1553 2018
rect 1598 2002 1601 2018
rect 1630 1992 1633 2018
rect 1646 2012 1649 2138
rect 1542 1960 1545 1979
rect 1574 1942 1577 1948
rect 1590 1932 1593 1938
rect 1510 1872 1513 1878
rect 1566 1872 1569 1908
rect 1606 1892 1609 1908
rect 1630 1902 1633 1988
rect 1662 1922 1665 2138
rect 1686 2132 1689 2138
rect 1710 2102 1713 2138
rect 1726 2132 1729 2138
rect 1758 2132 1761 2138
rect 1742 2122 1745 2128
rect 1710 2082 1713 2088
rect 1726 2062 1729 2068
rect 1758 2011 1761 2098
rect 1750 2008 1761 2011
rect 1750 1992 1753 2008
rect 1678 1952 1681 1988
rect 1718 1962 1721 1968
rect 1718 1942 1721 1948
rect 1734 1942 1737 1988
rect 1750 1958 1758 1961
rect 1742 1942 1745 1948
rect 1670 1912 1673 1918
rect 1642 1888 1646 1891
rect 1574 1882 1577 1888
rect 1614 1872 1617 1888
rect 1498 1868 1502 1871
rect 1550 1862 1553 1868
rect 1530 1858 1534 1861
rect 1494 1842 1497 1858
rect 1550 1842 1553 1848
rect 1566 1792 1569 1858
rect 1434 1768 1438 1771
rect 1510 1762 1513 1768
rect 1382 1742 1385 1748
rect 1326 1732 1329 1738
rect 1302 1682 1305 1688
rect 1310 1682 1313 1688
rect 1254 1672 1257 1678
rect 1278 1672 1281 1678
rect 1118 1652 1121 1658
rect 1062 1612 1065 1638
rect 1070 1572 1073 1578
rect 1046 1558 1054 1561
rect 1074 1558 1078 1561
rect 1094 1561 1097 1638
rect 1150 1632 1153 1658
rect 1102 1582 1105 1598
rect 1134 1592 1137 1618
rect 1110 1582 1113 1588
rect 1102 1572 1105 1578
rect 1166 1572 1169 1598
rect 1178 1588 1182 1591
rect 1198 1572 1201 1598
rect 1094 1558 1105 1561
rect 1030 1552 1033 1558
rect 1026 1548 1030 1551
rect 1006 1471 1009 1518
rect 1014 1502 1017 1518
rect 1006 1468 1014 1471
rect 1038 1462 1041 1538
rect 1046 1522 1049 1558
rect 1054 1552 1057 1558
rect 1086 1552 1089 1558
rect 1054 1492 1057 1538
rect 1062 1492 1065 1548
rect 1094 1541 1097 1548
rect 1086 1538 1097 1541
rect 1006 1442 1009 1458
rect 1038 1452 1041 1458
rect 1046 1452 1049 1488
rect 1070 1472 1073 1488
rect 1086 1472 1089 1538
rect 1054 1452 1057 1458
rect 1010 1438 1014 1441
rect 1026 1438 1030 1441
rect 1082 1418 1086 1421
rect 1006 1372 1009 1408
rect 1006 1352 1009 1368
rect 1038 1342 1041 1418
rect 1082 1358 1086 1361
rect 1046 1352 1049 1358
rect 1094 1352 1097 1518
rect 1102 1352 1105 1558
rect 1146 1558 1150 1561
rect 1118 1542 1121 1558
rect 1154 1548 1158 1551
rect 1126 1542 1129 1548
rect 1118 1442 1121 1538
rect 1138 1518 1142 1521
rect 1182 1492 1185 1558
rect 1190 1552 1193 1558
rect 1198 1512 1201 1518
rect 1206 1502 1209 1658
rect 1222 1562 1225 1668
rect 1242 1658 1246 1661
rect 1230 1642 1233 1648
rect 1238 1592 1241 1648
rect 1262 1642 1265 1648
rect 1278 1602 1281 1658
rect 1302 1632 1305 1678
rect 1270 1552 1273 1558
rect 1254 1542 1257 1548
rect 1266 1538 1273 1541
rect 1214 1532 1217 1538
rect 1270 1532 1273 1538
rect 1278 1532 1281 1558
rect 1286 1542 1289 1598
rect 1326 1582 1329 1728
rect 1338 1718 1342 1721
rect 1358 1711 1361 1738
rect 1366 1722 1369 1728
rect 1374 1712 1377 1718
rect 1390 1712 1393 1748
rect 1398 1722 1401 1748
rect 1414 1742 1417 1748
rect 1358 1708 1369 1711
rect 1338 1688 1342 1691
rect 1338 1658 1345 1661
rect 1298 1558 1302 1561
rect 1310 1552 1313 1558
rect 1294 1542 1297 1548
rect 1318 1542 1321 1578
rect 1222 1492 1225 1518
rect 1262 1492 1265 1528
rect 1126 1452 1129 1458
rect 1158 1362 1161 1418
rect 1150 1352 1153 1358
rect 1158 1352 1161 1358
rect 1058 1348 1062 1351
rect 1070 1342 1073 1348
rect 1094 1342 1097 1348
rect 1122 1338 1126 1341
rect 1022 1312 1025 1318
rect 966 1222 969 1238
rect 958 1158 969 1161
rect 902 1122 905 1138
rect 838 1072 841 1118
rect 862 1112 865 1118
rect 896 1103 898 1107
rect 902 1103 905 1107
rect 909 1103 912 1107
rect 854 1082 857 1088
rect 898 1058 902 1061
rect 790 1022 793 1048
rect 886 992 889 1008
rect 686 958 694 961
rect 702 932 705 938
rect 710 922 713 928
rect 678 872 681 878
rect 686 862 689 868
rect 674 858 678 861
rect 630 762 633 858
rect 686 822 689 848
rect 694 842 697 878
rect 710 852 713 908
rect 718 862 721 878
rect 622 702 625 748
rect 646 732 649 748
rect 654 712 657 738
rect 662 732 665 758
rect 670 742 673 748
rect 678 712 681 768
rect 698 748 702 751
rect 710 732 713 848
rect 726 842 729 978
rect 854 962 857 988
rect 894 962 897 1058
rect 918 1032 921 1148
rect 934 1092 937 1138
rect 942 1102 945 1158
rect 954 1148 958 1151
rect 954 1138 958 1141
rect 950 1122 953 1128
rect 942 992 945 1098
rect 966 1082 969 1158
rect 746 948 750 951
rect 806 942 809 948
rect 790 922 793 928
rect 758 872 761 878
rect 738 868 742 871
rect 774 862 777 898
rect 790 892 793 908
rect 802 878 806 881
rect 870 862 873 958
rect 902 942 905 948
rect 950 942 953 1078
rect 974 1071 977 1268
rect 1022 1232 1025 1308
rect 986 1148 990 1151
rect 1002 1148 1006 1151
rect 994 1138 998 1141
rect 982 1082 985 1118
rect 1006 1092 1009 1128
rect 1022 1112 1025 1118
rect 998 1082 1001 1088
rect 966 1068 977 1071
rect 1018 1068 1022 1071
rect 896 903 898 907
rect 902 903 905 907
rect 909 903 912 907
rect 926 872 929 878
rect 910 862 913 868
rect 754 858 758 861
rect 826 858 830 861
rect 762 848 766 851
rect 722 838 726 841
rect 722 818 726 821
rect 718 752 721 768
rect 726 762 729 788
rect 762 768 766 771
rect 774 762 777 858
rect 790 762 793 788
rect 746 748 750 751
rect 726 742 729 748
rect 718 732 721 738
rect 590 662 593 698
rect 630 682 633 688
rect 618 588 622 591
rect 630 582 633 678
rect 646 672 649 678
rect 694 622 697 648
rect 702 591 705 658
rect 710 652 713 728
rect 734 692 737 748
rect 766 732 769 738
rect 766 682 769 688
rect 774 682 777 758
rect 718 662 721 668
rect 750 662 753 668
rect 782 642 785 678
rect 782 592 785 638
rect 702 588 713 591
rect 710 552 713 588
rect 758 562 761 588
rect 790 552 793 618
rect 798 572 801 858
rect 806 662 809 858
rect 870 812 873 858
rect 878 831 881 850
rect 966 842 969 1068
rect 1006 1062 1009 1068
rect 986 1058 990 1061
rect 982 962 985 1018
rect 1014 1012 1017 1058
rect 974 952 977 958
rect 998 942 1001 998
rect 1022 982 1025 1058
rect 1030 1022 1033 1218
rect 1038 1212 1041 1338
rect 1054 1332 1057 1338
rect 1046 1262 1049 1268
rect 1038 1181 1041 1208
rect 1062 1182 1065 1218
rect 1038 1178 1049 1181
rect 1038 982 1041 1148
rect 1046 1142 1049 1178
rect 1070 1171 1073 1338
rect 1142 1332 1145 1338
rect 1086 1312 1089 1328
rect 1082 1288 1086 1291
rect 1102 1282 1105 1318
rect 1150 1292 1153 1338
rect 1166 1302 1169 1478
rect 1182 1421 1185 1468
rect 1214 1431 1217 1450
rect 1182 1418 1193 1421
rect 1182 1392 1185 1408
rect 1190 1402 1193 1418
rect 1206 1392 1209 1398
rect 1182 1352 1185 1388
rect 1190 1352 1193 1378
rect 1198 1342 1201 1378
rect 1194 1288 1198 1291
rect 1126 1272 1129 1278
rect 1182 1272 1185 1278
rect 1214 1272 1217 1398
rect 1254 1392 1257 1478
rect 1270 1472 1273 1528
rect 1286 1522 1289 1538
rect 1270 1432 1273 1468
rect 1278 1432 1281 1458
rect 1286 1452 1289 1458
rect 1222 1342 1225 1358
rect 1234 1348 1238 1351
rect 1230 1322 1233 1338
rect 1246 1322 1249 1358
rect 1258 1348 1262 1351
rect 1270 1342 1273 1388
rect 1294 1362 1297 1508
rect 1326 1492 1329 1548
rect 1334 1532 1337 1538
rect 1342 1512 1345 1658
rect 1350 1592 1353 1668
rect 1358 1652 1361 1658
rect 1366 1602 1369 1708
rect 1414 1682 1417 1688
rect 1382 1662 1385 1668
rect 1390 1652 1393 1668
rect 1398 1662 1401 1678
rect 1422 1672 1425 1698
rect 1446 1692 1449 1758
rect 1454 1752 1457 1758
rect 1482 1748 1494 1751
rect 1518 1732 1521 1758
rect 1534 1752 1537 1768
rect 1550 1752 1553 1778
rect 1582 1742 1585 1828
rect 1590 1802 1593 1858
rect 1610 1778 1614 1781
rect 1622 1752 1625 1858
rect 1630 1832 1633 1868
rect 1646 1862 1649 1878
rect 1654 1852 1657 1868
rect 1662 1862 1665 1898
rect 1678 1862 1681 1928
rect 1686 1872 1689 1878
rect 1670 1852 1673 1858
rect 1630 1792 1633 1808
rect 1610 1748 1614 1751
rect 1554 1738 1558 1741
rect 1526 1732 1529 1738
rect 1542 1732 1545 1738
rect 1562 1728 1566 1731
rect 1494 1702 1497 1718
rect 1494 1682 1497 1688
rect 1434 1678 1438 1681
rect 1542 1672 1545 1698
rect 1458 1668 1462 1671
rect 1470 1662 1473 1668
rect 1534 1662 1537 1668
rect 1550 1662 1553 1678
rect 1558 1672 1561 1718
rect 1590 1712 1593 1748
rect 1638 1742 1641 1848
rect 1694 1832 1697 1938
rect 1702 1872 1705 1908
rect 1710 1872 1713 1928
rect 1726 1881 1729 1918
rect 1726 1878 1737 1881
rect 1726 1862 1729 1868
rect 1702 1852 1705 1858
rect 1654 1792 1657 1798
rect 1718 1792 1721 1858
rect 1734 1842 1737 1878
rect 1742 1872 1745 1918
rect 1750 1882 1753 1958
rect 1746 1858 1750 1861
rect 1654 1752 1657 1778
rect 1734 1772 1737 1818
rect 1758 1812 1761 1938
rect 1766 1922 1769 2058
rect 1774 2022 1777 2048
rect 1782 2042 1785 2118
rect 1806 2082 1809 2118
rect 1838 2112 1841 2118
rect 1838 2072 1841 2088
rect 1846 2062 1849 2068
rect 1798 1972 1801 2018
rect 1806 1992 1809 2058
rect 1818 2048 1822 2051
rect 1830 2012 1833 2058
rect 1834 1988 1838 1991
rect 1774 1952 1777 1968
rect 1846 1952 1849 2008
rect 1782 1942 1785 1948
rect 1774 1892 1777 1898
rect 1766 1882 1769 1888
rect 1742 1772 1745 1778
rect 1782 1772 1785 1878
rect 1790 1802 1793 1948
rect 1798 1942 1801 1948
rect 1806 1932 1809 1938
rect 1798 1862 1801 1918
rect 1814 1912 1817 1918
rect 1854 1912 1857 2058
rect 1862 2012 1865 2148
rect 1950 2142 1953 2148
rect 1938 2138 1942 2141
rect 1986 2138 1990 2141
rect 2002 2138 2006 2141
rect 1878 2082 1881 2118
rect 1870 2062 1873 2068
rect 1870 2042 1873 2048
rect 1878 2042 1881 2068
rect 1886 2062 1889 2068
rect 1894 2062 1897 2138
rect 1918 2072 1921 2118
rect 1928 2103 1930 2107
rect 1934 2103 1937 2107
rect 1941 2103 1944 2107
rect 1902 2062 1905 2068
rect 1950 2062 1953 2098
rect 1958 2072 1961 2138
rect 2014 2132 2017 2158
rect 2022 2152 2025 2168
rect 2030 2141 2033 2218
rect 2054 2162 2057 2218
rect 2062 2202 2065 2328
rect 2086 2322 2089 2348
rect 2094 2332 2097 2468
rect 2118 2461 2121 2518
rect 2126 2502 2129 2548
rect 2134 2512 2137 2538
rect 2134 2492 2137 2508
rect 2142 2462 2145 2498
rect 2150 2481 2153 2538
rect 2166 2522 2169 2548
rect 2174 2542 2177 2558
rect 2158 2491 2161 2518
rect 2174 2502 2177 2528
rect 2174 2492 2177 2498
rect 2190 2492 2193 2638
rect 2198 2632 2201 2658
rect 2206 2652 2209 2658
rect 2214 2602 2217 2648
rect 2238 2601 2241 2618
rect 2238 2598 2246 2601
rect 2270 2592 2273 2658
rect 2294 2642 2297 2658
rect 2358 2652 2361 2668
rect 2382 2662 2385 2668
rect 2414 2662 2417 2668
rect 2326 2642 2329 2648
rect 2278 2622 2281 2628
rect 2322 2588 2326 2591
rect 2238 2552 2241 2588
rect 2334 2571 2337 2628
rect 2326 2568 2337 2571
rect 2342 2572 2345 2648
rect 2282 2558 2286 2561
rect 2282 2548 2286 2551
rect 2198 2532 2201 2548
rect 2218 2528 2222 2531
rect 2158 2488 2169 2491
rect 2166 2482 2169 2488
rect 2150 2478 2158 2481
rect 2114 2458 2121 2461
rect 2130 2458 2137 2461
rect 2110 2352 2113 2428
rect 2118 2372 2121 2418
rect 2126 2362 2129 2388
rect 2134 2352 2137 2458
rect 2142 2372 2145 2458
rect 2150 2362 2153 2478
rect 2222 2462 2225 2518
rect 2230 2492 2233 2548
rect 2318 2542 2321 2548
rect 2266 2528 2270 2531
rect 2254 2522 2257 2528
rect 2246 2481 2249 2518
rect 2262 2482 2265 2508
rect 2246 2478 2257 2481
rect 2246 2462 2249 2468
rect 2254 2462 2257 2478
rect 2262 2462 2265 2468
rect 2214 2452 2217 2458
rect 2158 2362 2161 2388
rect 2166 2352 2169 2428
rect 2222 2372 2225 2458
rect 2278 2392 2281 2538
rect 2302 2532 2305 2538
rect 2310 2532 2313 2538
rect 2310 2521 2313 2528
rect 2302 2518 2313 2521
rect 2294 2512 2297 2518
rect 2302 2492 2305 2518
rect 2310 2462 2313 2498
rect 2326 2472 2329 2568
rect 2334 2542 2337 2558
rect 2350 2552 2353 2598
rect 2366 2562 2369 2648
rect 2374 2632 2377 2658
rect 2422 2632 2425 2668
rect 2438 2662 2441 2748
rect 2430 2658 2438 2661
rect 2362 2548 2366 2551
rect 2398 2542 2401 2578
rect 2414 2562 2417 2608
rect 2422 2562 2425 2628
rect 2430 2592 2433 2658
rect 2454 2642 2457 2748
rect 2470 2731 2473 2748
rect 2478 2742 2481 2768
rect 2486 2742 2489 2838
rect 2494 2832 2497 2928
rect 2510 2902 2513 3078
rect 2526 3021 2529 3068
rect 2518 3018 2529 3021
rect 2558 3022 2561 3050
rect 2494 2792 2497 2828
rect 2506 2748 2510 2751
rect 2470 2728 2481 2731
rect 2478 2672 2481 2728
rect 2466 2668 2470 2671
rect 2440 2603 2442 2607
rect 2446 2603 2449 2607
rect 2453 2603 2456 2607
rect 2342 2532 2345 2538
rect 2426 2528 2430 2531
rect 2330 2458 2334 2461
rect 2318 2422 2321 2458
rect 2298 2418 2302 2421
rect 2174 2352 2177 2358
rect 2206 2352 2209 2368
rect 2238 2352 2241 2358
rect 2186 2348 2190 2351
rect 2226 2348 2230 2351
rect 2094 2282 2097 2298
rect 2102 2282 2105 2338
rect 2118 2282 2121 2348
rect 2130 2338 2134 2341
rect 2142 2312 2145 2348
rect 2078 2262 2081 2278
rect 2102 2262 2105 2278
rect 2142 2262 2145 2308
rect 2182 2301 2185 2338
rect 2174 2298 2185 2301
rect 2137 2258 2142 2261
rect 2074 2248 2078 2251
rect 2042 2158 2046 2161
rect 2042 2148 2046 2151
rect 2030 2138 2038 2141
rect 2050 2138 2054 2141
rect 1966 2061 1969 2078
rect 1978 2068 1982 2071
rect 1958 2058 1969 2061
rect 1990 2062 1993 2098
rect 1938 2048 1942 2051
rect 1886 2011 1889 2018
rect 1886 2008 1894 2011
rect 1866 1988 1870 1991
rect 1878 1952 1881 2008
rect 1950 1961 1953 2018
rect 1946 1958 1953 1961
rect 1958 1992 1961 2058
rect 2006 2042 2009 2078
rect 2014 2052 2017 2068
rect 2022 2062 2025 2098
rect 2038 2062 2041 2068
rect 1994 2038 1998 2041
rect 2038 2041 2041 2048
rect 2030 2038 2041 2041
rect 1966 1992 1969 1998
rect 1930 1948 1934 1951
rect 1906 1938 1910 1941
rect 1958 1932 1961 1988
rect 1974 1932 1977 1978
rect 1982 1962 1985 1968
rect 1998 1942 2001 1958
rect 2006 1952 2009 2038
rect 2030 2011 2033 2038
rect 2046 2012 2049 2078
rect 2054 2052 2057 2128
rect 2062 2102 2065 2148
rect 2070 2142 2073 2168
rect 2078 2142 2081 2168
rect 2086 2141 2089 2218
rect 2094 2172 2097 2228
rect 2126 2152 2129 2258
rect 2110 2142 2113 2148
rect 2086 2138 2094 2141
rect 2122 2138 2126 2141
rect 2090 2128 2094 2131
rect 2082 2088 2086 2091
rect 2126 2082 2129 2118
rect 2102 2078 2110 2081
rect 2078 2062 2081 2068
rect 2102 2062 2105 2078
rect 2114 2068 2118 2071
rect 2126 2062 2129 2068
rect 2066 2058 2070 2061
rect 2030 2008 2038 2011
rect 2014 1952 2017 1958
rect 1994 1938 1998 1941
rect 2014 1932 2017 1938
rect 2030 1922 2033 2008
rect 2038 1942 2041 1948
rect 2046 1942 2049 2008
rect 2054 1992 2057 2048
rect 2070 1952 2073 1998
rect 1946 1918 1953 1921
rect 1894 1902 1897 1918
rect 1928 1903 1930 1907
rect 1934 1903 1937 1907
rect 1941 1903 1944 1907
rect 1870 1882 1873 1888
rect 1854 1852 1857 1868
rect 1910 1862 1913 1888
rect 1822 1831 1825 1850
rect 1774 1762 1777 1768
rect 1598 1722 1601 1728
rect 1646 1702 1649 1738
rect 1566 1662 1569 1688
rect 1578 1678 1582 1681
rect 1406 1658 1414 1661
rect 1434 1658 1438 1661
rect 1482 1658 1486 1661
rect 1506 1658 1510 1661
rect 1358 1542 1361 1578
rect 1374 1551 1377 1638
rect 1370 1548 1377 1551
rect 1390 1542 1393 1598
rect 1406 1591 1409 1658
rect 1416 1603 1418 1607
rect 1422 1603 1425 1607
rect 1429 1603 1432 1607
rect 1406 1588 1414 1591
rect 1354 1528 1358 1531
rect 1366 1522 1369 1528
rect 1390 1512 1393 1538
rect 1342 1492 1345 1498
rect 1294 1352 1297 1358
rect 1302 1352 1305 1418
rect 1310 1361 1313 1478
rect 1350 1472 1353 1498
rect 1366 1492 1369 1508
rect 1398 1482 1401 1488
rect 1414 1482 1417 1528
rect 1430 1492 1433 1558
rect 1454 1552 1457 1598
rect 1446 1532 1449 1538
rect 1438 1522 1441 1528
rect 1358 1472 1361 1478
rect 1318 1452 1321 1468
rect 1362 1458 1366 1461
rect 1318 1402 1321 1448
rect 1326 1392 1329 1458
rect 1342 1392 1345 1458
rect 1382 1442 1385 1458
rect 1390 1452 1393 1468
rect 1310 1358 1318 1361
rect 1342 1352 1345 1358
rect 1350 1352 1353 1358
rect 1374 1352 1377 1408
rect 1390 1392 1393 1448
rect 1406 1412 1409 1448
rect 1422 1442 1425 1478
rect 1446 1472 1449 1508
rect 1454 1461 1457 1548
rect 1462 1492 1465 1658
rect 1470 1562 1473 1598
rect 1478 1572 1481 1658
rect 1482 1538 1486 1541
rect 1470 1502 1473 1518
rect 1502 1492 1505 1648
rect 1574 1612 1577 1668
rect 1590 1651 1593 1678
rect 1598 1672 1601 1698
rect 1622 1662 1625 1688
rect 1630 1672 1633 1678
rect 1654 1662 1657 1708
rect 1670 1692 1673 1748
rect 1678 1742 1681 1758
rect 1726 1752 1729 1758
rect 1686 1742 1689 1748
rect 1706 1738 1710 1741
rect 1734 1732 1737 1758
rect 1778 1748 1782 1751
rect 1698 1728 1702 1731
rect 1662 1672 1665 1678
rect 1670 1672 1673 1688
rect 1710 1672 1713 1728
rect 1726 1682 1729 1688
rect 1734 1681 1737 1728
rect 1750 1692 1753 1728
rect 1734 1678 1742 1681
rect 1758 1681 1761 1738
rect 1814 1722 1817 1798
rect 1918 1752 1921 1888
rect 1950 1872 1953 1918
rect 1958 1832 1961 1858
rect 1934 1762 1937 1788
rect 1886 1732 1889 1738
rect 1870 1722 1873 1728
rect 1786 1718 1790 1721
rect 1750 1678 1761 1681
rect 1610 1658 1614 1661
rect 1630 1658 1638 1661
rect 1590 1648 1601 1651
rect 1610 1648 1614 1651
rect 1566 1592 1569 1598
rect 1510 1552 1513 1558
rect 1518 1552 1521 1588
rect 1530 1568 1534 1571
rect 1542 1552 1545 1558
rect 1566 1552 1569 1568
rect 1582 1562 1585 1568
rect 1590 1552 1593 1638
rect 1598 1632 1601 1648
rect 1622 1592 1625 1608
rect 1602 1568 1606 1571
rect 1614 1562 1617 1568
rect 1554 1548 1558 1551
rect 1630 1542 1633 1658
rect 1638 1612 1641 1648
rect 1638 1562 1641 1608
rect 1554 1538 1558 1541
rect 1590 1532 1593 1538
rect 1474 1488 1478 1491
rect 1486 1482 1489 1488
rect 1530 1478 1534 1481
rect 1614 1472 1617 1538
rect 1630 1481 1633 1528
rect 1638 1512 1641 1518
rect 1646 1492 1649 1648
rect 1654 1542 1657 1548
rect 1662 1542 1665 1668
rect 1710 1642 1713 1658
rect 1670 1502 1673 1638
rect 1718 1632 1721 1668
rect 1678 1572 1681 1618
rect 1694 1562 1697 1608
rect 1678 1552 1681 1558
rect 1686 1502 1689 1538
rect 1686 1482 1689 1488
rect 1702 1482 1705 1538
rect 1710 1512 1713 1548
rect 1626 1478 1633 1481
rect 1670 1472 1673 1478
rect 1710 1472 1713 1488
rect 1718 1482 1721 1628
rect 1726 1552 1729 1558
rect 1734 1552 1737 1658
rect 1750 1652 1753 1678
rect 1758 1562 1761 1658
rect 1774 1632 1777 1638
rect 1774 1612 1777 1628
rect 1774 1562 1777 1568
rect 1750 1552 1753 1558
rect 1746 1538 1750 1541
rect 1734 1502 1737 1538
rect 1766 1492 1769 1518
rect 1754 1478 1758 1481
rect 1498 1468 1502 1471
rect 1578 1468 1582 1471
rect 1682 1468 1686 1471
rect 1454 1458 1465 1461
rect 1450 1448 1454 1451
rect 1416 1403 1418 1407
rect 1422 1403 1425 1407
rect 1429 1403 1432 1407
rect 1298 1338 1302 1341
rect 1230 1282 1233 1288
rect 1270 1272 1273 1338
rect 1278 1272 1281 1318
rect 1286 1272 1289 1278
rect 1094 1252 1097 1268
rect 1078 1242 1081 1248
rect 1102 1222 1105 1268
rect 1158 1262 1161 1268
rect 1190 1262 1193 1268
rect 1262 1262 1265 1268
rect 1294 1262 1297 1318
rect 1310 1272 1313 1318
rect 1318 1272 1321 1348
rect 1130 1258 1134 1261
rect 1206 1252 1209 1258
rect 1178 1248 1182 1251
rect 1110 1182 1113 1218
rect 1070 1168 1081 1171
rect 1070 1152 1073 1158
rect 1078 1152 1081 1168
rect 1118 1162 1121 1248
rect 1150 1242 1153 1248
rect 1162 1238 1166 1241
rect 1246 1222 1249 1258
rect 1098 1158 1102 1161
rect 1058 1148 1062 1151
rect 1122 1148 1126 1151
rect 1078 1142 1081 1148
rect 1110 1142 1113 1148
rect 1134 1141 1137 1208
rect 1142 1152 1145 1158
rect 1134 1138 1142 1141
rect 1086 1132 1089 1138
rect 1102 1132 1105 1138
rect 1046 1062 1049 1068
rect 1054 1062 1057 1118
rect 1070 1082 1073 1118
rect 1110 1062 1113 1108
rect 1058 1048 1062 1051
rect 1050 1028 1054 1031
rect 1070 1012 1073 1058
rect 1078 1042 1081 1048
rect 1054 992 1057 1008
rect 1022 962 1025 968
rect 1030 952 1033 978
rect 1006 942 1009 948
rect 974 852 977 918
rect 982 882 985 918
rect 1006 892 1009 928
rect 1018 918 1022 921
rect 1018 878 1022 881
rect 894 752 897 808
rect 838 732 841 738
rect 854 722 857 728
rect 878 692 881 708
rect 896 703 898 707
rect 902 703 905 707
rect 909 703 912 707
rect 926 692 929 818
rect 934 792 937 798
rect 818 668 822 671
rect 838 662 841 668
rect 886 662 889 678
rect 934 662 937 778
rect 966 742 969 838
rect 958 682 961 688
rect 822 652 825 658
rect 834 648 838 651
rect 854 641 857 658
rect 850 638 857 641
rect 838 592 841 618
rect 854 592 857 638
rect 806 562 809 588
rect 814 562 817 568
rect 862 552 865 658
rect 870 552 873 558
rect 842 548 846 551
rect 542 538 553 541
rect 570 538 574 541
rect 486 392 489 408
rect 526 392 529 418
rect 534 392 537 538
rect 542 462 545 538
rect 562 438 566 441
rect 386 268 390 271
rect 410 258 414 261
rect 346 218 350 221
rect 314 188 318 191
rect 182 160 185 179
rect 142 132 145 138
rect 142 82 145 128
rect 166 102 169 148
rect 214 142 217 148
rect 230 122 233 128
rect 30 72 33 78
rect 158 72 161 78
rect 198 62 201 98
rect 230 62 233 108
rect 310 92 313 178
rect 342 152 345 158
rect 254 72 257 78
rect 6 42 9 48
rect 190 22 193 50
rect 326 32 329 118
rect 350 82 353 118
rect 342 62 345 68
rect 358 61 361 228
rect 374 72 377 218
rect 392 203 394 207
rect 398 203 401 207
rect 405 203 408 207
rect 414 62 417 208
rect 354 58 361 61
rect 378 58 382 61
rect 238 -19 242 -18
rect 246 -19 249 18
rect 238 -22 249 -19
rect 326 -18 329 18
rect 342 -18 345 28
rect 410 18 417 21
rect 358 -18 361 8
rect 326 -22 330 -18
rect 342 -22 346 -18
rect 358 -22 362 -18
rect 366 -19 369 18
rect 392 3 394 7
rect 398 3 401 7
rect 405 3 408 7
rect 414 -18 417 18
rect 374 -19 378 -18
rect 366 -22 378 -19
rect 414 -22 418 -18
rect 422 -19 425 218
rect 438 212 441 218
rect 478 132 481 388
rect 558 362 561 428
rect 574 402 577 418
rect 582 352 585 548
rect 522 348 526 351
rect 590 342 593 538
rect 710 532 713 538
rect 694 522 697 528
rect 598 352 601 518
rect 694 502 697 518
rect 654 482 657 488
rect 742 472 745 548
rect 802 538 806 541
rect 834 538 838 541
rect 782 522 785 538
rect 670 442 673 468
rect 718 462 721 468
rect 738 458 742 461
rect 702 422 705 450
rect 614 362 617 398
rect 646 352 649 358
rect 678 352 681 358
rect 618 348 622 351
rect 530 338 534 341
rect 502 322 505 328
rect 534 292 537 318
rect 518 282 521 288
rect 534 272 537 278
rect 582 262 585 298
rect 526 160 529 179
rect 534 152 537 258
rect 566 231 569 250
rect 582 152 585 258
rect 614 232 617 318
rect 630 262 633 298
rect 638 272 641 318
rect 662 302 665 318
rect 686 282 689 388
rect 694 332 697 338
rect 722 318 726 321
rect 670 272 673 278
rect 686 252 689 278
rect 638 231 641 250
rect 494 142 497 148
rect 566 102 569 118
rect 526 82 529 88
rect 542 62 545 68
rect 582 62 585 148
rect 614 122 617 218
rect 634 148 638 151
rect 678 132 681 208
rect 726 160 729 179
rect 694 142 697 148
rect 442 58 445 61
rect 614 52 617 118
rect 638 82 641 108
rect 638 72 641 78
rect 734 72 737 168
rect 750 82 753 498
rect 758 492 761 518
rect 782 402 785 418
rect 758 302 761 348
rect 798 332 801 418
rect 814 382 817 518
rect 886 502 889 518
rect 896 503 898 507
rect 902 503 905 507
rect 909 503 912 507
rect 862 482 865 488
rect 822 402 825 458
rect 878 422 881 468
rect 910 431 913 450
rect 846 352 849 398
rect 862 362 865 388
rect 894 372 897 378
rect 926 362 929 648
rect 934 612 937 658
rect 934 562 937 588
rect 898 348 902 351
rect 814 342 817 348
rect 846 322 849 348
rect 886 342 889 348
rect 926 342 929 358
rect 770 288 774 291
rect 782 262 785 298
rect 838 282 841 288
rect 854 282 857 328
rect 896 303 898 307
rect 902 303 905 307
rect 909 303 912 307
rect 806 272 809 278
rect 818 268 822 271
rect 790 192 793 198
rect 790 162 793 188
rect 766 102 769 118
rect 630 62 633 68
rect 682 58 686 61
rect 574 31 577 50
rect 638 51 641 58
rect 634 48 641 51
rect 702 31 705 50
rect 430 12 433 18
rect 446 -18 449 8
rect 542 -18 545 8
rect 558 -18 561 8
rect 574 -18 577 8
rect 630 -18 633 8
rect 430 -19 434 -18
rect 422 -22 434 -19
rect 446 -22 450 -18
rect 542 -22 546 -18
rect 558 -22 562 -18
rect 574 -22 578 -18
rect 630 -22 634 -18
rect 654 -19 658 -18
rect 662 -19 665 18
rect 654 -22 665 -19
rect 774 -18 777 8
rect 774 -22 778 -18
rect 790 -19 794 -18
rect 798 -19 801 218
rect 806 162 809 268
rect 830 262 833 268
rect 818 258 822 261
rect 830 232 833 248
rect 830 172 833 178
rect 806 72 809 148
rect 822 142 825 158
rect 830 142 833 148
rect 814 112 817 138
rect 838 131 841 278
rect 854 272 857 278
rect 922 268 926 271
rect 854 222 857 268
rect 866 258 873 261
rect 898 258 902 261
rect 862 242 865 248
rect 870 192 873 258
rect 878 212 881 248
rect 846 162 849 168
rect 886 162 889 248
rect 894 232 897 238
rect 902 212 905 238
rect 894 192 897 208
rect 902 172 905 208
rect 934 192 937 488
rect 950 402 953 658
rect 966 602 969 738
rect 998 672 1001 718
rect 974 662 977 668
rect 982 642 985 668
rect 1006 662 1009 798
rect 1022 792 1025 868
rect 1030 832 1033 938
rect 1046 882 1049 988
rect 1058 948 1062 951
rect 1070 942 1073 948
rect 1038 852 1041 858
rect 1038 762 1041 818
rect 1062 812 1065 938
rect 1070 932 1073 938
rect 1078 742 1081 938
rect 1086 912 1089 1018
rect 1094 992 1097 998
rect 1094 932 1097 938
rect 1102 901 1105 1058
rect 1110 1022 1113 1048
rect 1110 952 1113 958
rect 1118 912 1121 1118
rect 1158 1072 1161 1208
rect 1166 1152 1169 1218
rect 1182 1160 1185 1179
rect 1166 1112 1169 1148
rect 1278 1142 1281 1258
rect 1214 1132 1217 1138
rect 1294 1132 1297 1218
rect 1302 1152 1305 1268
rect 1310 1232 1313 1248
rect 1310 1192 1313 1198
rect 1230 1122 1233 1128
rect 1254 1092 1257 1108
rect 1174 1042 1177 1078
rect 1270 1062 1273 1068
rect 1278 1062 1281 1078
rect 1302 1071 1305 1148
rect 1318 1142 1321 1268
rect 1326 1262 1329 1318
rect 1326 1162 1329 1218
rect 1334 1192 1337 1328
rect 1342 1292 1345 1348
rect 1374 1341 1377 1348
rect 1370 1338 1377 1341
rect 1390 1342 1393 1378
rect 1414 1362 1417 1378
rect 1426 1358 1430 1361
rect 1394 1338 1398 1341
rect 1390 1292 1393 1298
rect 1362 1288 1366 1291
rect 1350 1272 1353 1278
rect 1366 1272 1369 1278
rect 1398 1272 1401 1278
rect 1342 1252 1345 1268
rect 1374 1262 1377 1268
rect 1402 1258 1406 1261
rect 1358 1192 1361 1248
rect 1334 1152 1337 1158
rect 1302 1068 1310 1071
rect 1298 1058 1302 1061
rect 1302 1052 1305 1058
rect 1142 952 1145 998
rect 1174 962 1177 998
rect 1198 952 1201 958
rect 1214 952 1217 988
rect 1222 952 1225 958
rect 1130 948 1134 951
rect 1154 948 1158 951
rect 1186 948 1190 951
rect 1250 948 1254 951
rect 1266 948 1270 951
rect 1142 942 1145 948
rect 1234 938 1238 941
rect 1126 932 1129 938
rect 1150 932 1153 938
rect 1166 922 1169 938
rect 1094 898 1105 901
rect 1094 862 1097 898
rect 1134 882 1137 888
rect 1150 872 1153 878
rect 1222 872 1225 938
rect 1262 932 1265 938
rect 1230 892 1233 918
rect 1262 872 1265 918
rect 1278 892 1281 1048
rect 1310 1042 1313 1068
rect 1294 961 1297 1018
rect 1294 958 1305 961
rect 1286 952 1289 958
rect 1302 952 1305 958
rect 1294 942 1297 948
rect 1294 932 1297 938
rect 1286 882 1289 918
rect 1294 872 1297 878
rect 1182 822 1185 850
rect 1102 792 1105 808
rect 1206 782 1209 858
rect 1194 768 1198 771
rect 1174 762 1177 768
rect 1210 758 1214 761
rect 1078 732 1081 738
rect 1066 728 1070 731
rect 1038 702 1041 718
rect 1078 692 1081 728
rect 1086 702 1089 748
rect 1118 742 1121 748
rect 1126 732 1129 758
rect 1142 732 1145 738
rect 1150 722 1153 748
rect 1158 742 1161 758
rect 1174 742 1177 748
rect 1106 718 1110 721
rect 1134 702 1137 718
rect 1110 672 1113 678
rect 1126 672 1129 678
rect 1026 658 1030 661
rect 998 652 1001 658
rect 1038 652 1041 658
rect 1026 638 1030 641
rect 1078 631 1081 650
rect 1014 622 1017 628
rect 1082 588 1086 591
rect 982 542 985 568
rect 998 532 1001 578
rect 1090 558 1094 561
rect 1110 552 1113 658
rect 1042 548 1046 551
rect 1118 542 1121 618
rect 1126 562 1129 668
rect 1166 662 1169 718
rect 1198 702 1201 748
rect 1222 742 1225 828
rect 1218 738 1221 741
rect 1238 712 1241 838
rect 1246 732 1249 848
rect 1270 822 1273 868
rect 1302 862 1305 888
rect 1310 882 1313 1038
rect 1318 962 1321 1108
rect 1326 1062 1329 1078
rect 1334 1062 1337 1068
rect 1342 1062 1345 1168
rect 1350 1162 1353 1168
rect 1374 1162 1377 1258
rect 1394 1248 1398 1251
rect 1414 1221 1417 1318
rect 1422 1252 1425 1328
rect 1438 1282 1441 1438
rect 1446 1332 1449 1358
rect 1462 1352 1465 1458
rect 1454 1342 1457 1348
rect 1462 1322 1465 1348
rect 1470 1312 1473 1468
rect 1514 1458 1518 1461
rect 1526 1451 1529 1468
rect 1598 1462 1601 1468
rect 1570 1458 1574 1461
rect 1586 1458 1590 1461
rect 1658 1458 1662 1461
rect 1678 1458 1686 1461
rect 1746 1458 1750 1461
rect 1518 1448 1529 1451
rect 1510 1442 1513 1448
rect 1502 1382 1505 1388
rect 1478 1362 1481 1378
rect 1482 1348 1486 1351
rect 1482 1318 1486 1321
rect 1446 1278 1473 1281
rect 1446 1272 1449 1278
rect 1470 1271 1473 1278
rect 1470 1268 1478 1271
rect 1498 1268 1502 1271
rect 1462 1262 1465 1268
rect 1510 1262 1513 1268
rect 1458 1258 1462 1261
rect 1474 1258 1478 1261
rect 1490 1248 1494 1251
rect 1406 1218 1417 1221
rect 1406 1212 1409 1218
rect 1416 1203 1418 1207
rect 1422 1203 1425 1207
rect 1429 1203 1432 1207
rect 1438 1172 1441 1178
rect 1422 1152 1425 1158
rect 1494 1152 1497 1198
rect 1502 1192 1505 1258
rect 1510 1232 1513 1248
rect 1510 1192 1513 1228
rect 1518 1192 1521 1448
rect 1558 1392 1561 1408
rect 1526 1302 1529 1348
rect 1550 1342 1553 1358
rect 1542 1312 1545 1318
rect 1534 1282 1537 1298
rect 1534 1272 1537 1278
rect 1526 1262 1529 1268
rect 1542 1252 1545 1268
rect 1550 1252 1553 1258
rect 1558 1241 1561 1378
rect 1574 1342 1577 1408
rect 1638 1402 1641 1458
rect 1650 1448 1654 1451
rect 1590 1352 1593 1398
rect 1606 1352 1609 1388
rect 1574 1332 1577 1338
rect 1566 1322 1569 1328
rect 1574 1272 1577 1308
rect 1590 1281 1593 1348
rect 1610 1318 1614 1321
rect 1582 1278 1593 1281
rect 1566 1262 1569 1268
rect 1582 1262 1585 1278
rect 1550 1238 1561 1241
rect 1566 1242 1569 1248
rect 1550 1192 1553 1238
rect 1566 1202 1569 1238
rect 1458 1148 1462 1151
rect 1350 1112 1353 1118
rect 1358 1092 1361 1108
rect 1350 1072 1353 1088
rect 1366 1082 1369 1128
rect 1374 1072 1377 1118
rect 1382 1112 1385 1118
rect 1402 1088 1406 1091
rect 1422 1082 1425 1108
rect 1382 1062 1385 1068
rect 1342 982 1345 1058
rect 1390 1052 1393 1078
rect 1430 1062 1433 1098
rect 1446 1092 1449 1148
rect 1458 1138 1462 1141
rect 1482 1138 1486 1141
rect 1498 1128 1502 1131
rect 1474 1118 1478 1121
rect 1438 1062 1441 1068
rect 1354 1048 1358 1051
rect 1326 962 1329 968
rect 1358 952 1361 958
rect 1374 952 1377 998
rect 1390 952 1393 1008
rect 1406 992 1409 1058
rect 1416 1003 1418 1007
rect 1422 1003 1425 1007
rect 1429 1003 1432 1007
rect 1446 962 1449 1088
rect 1462 1062 1465 1098
rect 1474 1068 1478 1071
rect 1502 1062 1505 1118
rect 1510 1092 1513 1118
rect 1518 1102 1521 1148
rect 1542 1132 1545 1138
rect 1530 1128 1534 1131
rect 1550 1102 1553 1148
rect 1566 1132 1569 1158
rect 1574 1152 1577 1178
rect 1582 1162 1585 1218
rect 1598 1172 1601 1248
rect 1606 1212 1609 1278
rect 1622 1272 1625 1358
rect 1630 1342 1633 1348
rect 1638 1322 1641 1328
rect 1646 1272 1649 1358
rect 1654 1352 1657 1398
rect 1654 1262 1657 1268
rect 1626 1258 1630 1261
rect 1614 1192 1617 1248
rect 1638 1241 1641 1258
rect 1626 1238 1641 1241
rect 1590 1122 1593 1128
rect 1606 1122 1609 1138
rect 1518 1062 1521 1098
rect 1570 1088 1574 1091
rect 1534 1082 1537 1088
rect 1550 1072 1553 1088
rect 1574 1072 1577 1078
rect 1538 1068 1542 1071
rect 1482 1058 1486 1061
rect 1526 1061 1529 1068
rect 1582 1062 1585 1118
rect 1614 1102 1617 1148
rect 1622 1092 1625 1218
rect 1630 1132 1633 1158
rect 1638 1142 1641 1198
rect 1662 1192 1665 1358
rect 1670 1352 1673 1388
rect 1678 1291 1681 1458
rect 1686 1352 1689 1428
rect 1702 1392 1705 1438
rect 1718 1362 1721 1378
rect 1694 1342 1697 1348
rect 1686 1302 1689 1338
rect 1694 1318 1702 1321
rect 1678 1288 1689 1291
rect 1670 1202 1673 1258
rect 1678 1192 1681 1238
rect 1638 1092 1641 1138
rect 1646 1122 1649 1148
rect 1526 1058 1534 1061
rect 1470 1022 1473 1058
rect 1510 1051 1513 1058
rect 1606 1052 1609 1068
rect 1622 1052 1625 1078
rect 1646 1072 1649 1078
rect 1506 1048 1513 1051
rect 1570 1048 1582 1051
rect 1534 992 1537 1008
rect 1498 958 1502 961
rect 1446 952 1449 958
rect 1342 932 1345 948
rect 1350 942 1353 948
rect 1318 902 1321 918
rect 1326 902 1329 918
rect 1330 888 1334 891
rect 1342 882 1345 888
rect 1350 872 1353 878
rect 1358 872 1361 948
rect 1366 922 1369 948
rect 1434 938 1438 941
rect 1378 928 1382 931
rect 1406 882 1409 888
rect 1430 882 1433 928
rect 1454 912 1457 938
rect 1462 922 1465 958
rect 1478 952 1481 958
rect 1490 948 1494 951
rect 1474 938 1478 941
rect 1458 888 1465 891
rect 1462 882 1465 888
rect 1314 858 1318 861
rect 1306 838 1310 841
rect 1254 762 1257 818
rect 1286 812 1289 838
rect 1326 792 1329 868
rect 1370 858 1374 861
rect 1350 802 1353 858
rect 1362 848 1366 851
rect 1382 841 1385 868
rect 1390 852 1393 858
rect 1382 838 1393 841
rect 1262 752 1265 778
rect 1350 760 1353 779
rect 1374 752 1377 838
rect 1390 792 1393 838
rect 1430 822 1433 878
rect 1458 868 1462 871
rect 1478 862 1481 928
rect 1458 858 1462 861
rect 1416 803 1418 807
rect 1422 803 1425 807
rect 1429 803 1432 807
rect 1406 792 1409 798
rect 1426 788 1430 791
rect 1470 752 1473 768
rect 1478 762 1481 858
rect 1486 812 1489 938
rect 1510 932 1513 938
rect 1526 932 1529 948
rect 1494 892 1497 908
rect 1494 842 1497 858
rect 1486 752 1489 808
rect 1502 792 1505 888
rect 1510 862 1513 868
rect 1526 852 1529 898
rect 1458 748 1462 751
rect 1302 732 1305 748
rect 1494 742 1497 758
rect 1466 738 1470 741
rect 1482 738 1486 741
rect 1318 732 1321 738
rect 1238 692 1241 698
rect 1246 692 1249 728
rect 1242 668 1246 671
rect 1282 668 1286 671
rect 1214 652 1217 658
rect 1230 652 1233 668
rect 1254 651 1257 658
rect 1250 648 1257 651
rect 1262 652 1265 658
rect 1270 632 1273 668
rect 1294 662 1297 698
rect 1314 658 1318 661
rect 1286 652 1289 658
rect 1334 652 1337 688
rect 1350 672 1353 738
rect 1494 732 1497 738
rect 1374 672 1377 678
rect 1310 642 1313 648
rect 1202 618 1206 621
rect 1142 552 1145 598
rect 1182 560 1185 579
rect 1158 552 1161 558
rect 1274 548 1278 551
rect 974 482 977 508
rect 982 472 985 518
rect 990 462 993 478
rect 950 372 953 398
rect 942 352 945 358
rect 966 352 969 418
rect 974 362 977 368
rect 982 351 985 458
rect 1014 452 1017 488
rect 1046 482 1049 488
rect 1022 452 1025 458
rect 990 442 993 448
rect 1054 442 1057 478
rect 1070 442 1073 498
rect 1078 462 1081 488
rect 1086 452 1089 528
rect 1126 522 1129 528
rect 1114 488 1118 491
rect 1126 472 1129 518
rect 1142 492 1145 548
rect 1134 472 1137 478
rect 1166 472 1169 518
rect 1214 482 1217 538
rect 1230 532 1233 538
rect 1302 522 1305 618
rect 1310 582 1313 588
rect 1326 552 1329 558
rect 1334 552 1337 618
rect 1350 592 1353 658
rect 1358 582 1361 668
rect 1382 652 1385 678
rect 1390 662 1393 708
rect 1398 702 1401 728
rect 1430 712 1433 728
rect 1446 692 1449 728
rect 1442 678 1454 681
rect 1450 668 1454 671
rect 1430 662 1433 668
rect 1462 662 1465 728
rect 1502 712 1505 748
rect 1494 682 1497 708
rect 1470 672 1473 678
rect 1486 672 1489 678
rect 1270 482 1273 488
rect 1254 472 1257 478
rect 978 348 985 351
rect 966 342 969 348
rect 998 342 1001 378
rect 1014 362 1017 418
rect 1030 402 1033 438
rect 1062 412 1065 418
rect 1094 402 1097 458
rect 1102 442 1105 468
rect 1070 362 1073 368
rect 1042 358 1046 361
rect 982 262 985 318
rect 1014 302 1017 358
rect 1026 348 1030 351
rect 1054 342 1057 358
rect 1062 342 1065 348
rect 1086 332 1089 338
rect 1046 272 1049 278
rect 1030 262 1033 268
rect 1086 262 1089 318
rect 1094 302 1097 358
rect 1110 342 1113 468
rect 1142 462 1145 468
rect 1166 462 1169 468
rect 1134 451 1137 458
rect 1182 452 1185 468
rect 1130 448 1137 451
rect 1142 442 1145 448
rect 1130 388 1134 391
rect 1190 372 1193 378
rect 1142 362 1145 368
rect 1182 352 1185 358
rect 1190 352 1193 358
rect 1198 352 1201 368
rect 1146 348 1150 351
rect 954 258 958 261
rect 934 162 937 188
rect 942 182 945 258
rect 962 248 966 251
rect 998 231 1001 250
rect 950 172 953 208
rect 962 168 966 171
rect 1010 168 1014 171
rect 890 158 894 161
rect 978 158 982 161
rect 942 152 945 158
rect 850 148 854 151
rect 898 148 902 151
rect 978 148 982 151
rect 990 142 993 158
rect 1010 148 1014 151
rect 1022 142 1025 158
rect 1030 142 1033 218
rect 1038 162 1041 168
rect 1054 162 1057 168
rect 1038 142 1041 148
rect 962 138 966 141
rect 998 132 1001 138
rect 1062 132 1065 198
rect 1086 192 1089 258
rect 1094 212 1097 298
rect 1118 282 1121 348
rect 1126 342 1129 348
rect 1150 282 1153 328
rect 1134 272 1137 278
rect 1166 271 1169 318
rect 1198 302 1201 348
rect 1214 322 1217 458
rect 1310 452 1313 518
rect 1222 431 1225 450
rect 1222 332 1225 408
rect 1238 362 1241 368
rect 1286 362 1289 368
rect 1230 342 1233 348
rect 1238 322 1241 348
rect 1254 292 1257 358
rect 1262 352 1265 358
rect 1294 352 1297 408
rect 1326 382 1329 548
rect 1358 472 1361 548
rect 1374 542 1377 578
rect 1382 572 1385 578
rect 1390 572 1393 658
rect 1422 642 1425 658
rect 1422 622 1425 638
rect 1406 552 1409 618
rect 1416 603 1418 607
rect 1422 603 1425 607
rect 1429 603 1432 607
rect 1438 602 1441 658
rect 1414 552 1417 558
rect 1386 548 1390 551
rect 1438 551 1441 598
rect 1446 562 1449 568
rect 1434 548 1441 551
rect 1454 552 1457 658
rect 1478 652 1481 668
rect 1494 662 1497 668
rect 1462 592 1465 648
rect 1486 592 1489 638
rect 1482 548 1486 551
rect 1426 538 1430 541
rect 1374 532 1377 538
rect 1398 472 1401 528
rect 1414 472 1417 478
rect 1386 458 1390 461
rect 1314 368 1318 371
rect 1334 362 1337 448
rect 1354 418 1358 421
rect 1374 372 1377 418
rect 1350 362 1353 368
rect 1318 352 1321 358
rect 1334 342 1337 358
rect 1350 342 1353 348
rect 1270 302 1273 338
rect 1286 332 1289 338
rect 1306 328 1310 331
rect 1158 268 1169 271
rect 1174 272 1177 278
rect 1230 272 1233 278
rect 1290 268 1294 271
rect 1078 162 1081 188
rect 1086 172 1089 178
rect 1094 172 1097 208
rect 1110 172 1113 218
rect 1118 192 1121 258
rect 1158 232 1161 268
rect 1166 242 1169 258
rect 1182 252 1185 268
rect 1206 262 1209 268
rect 1214 262 1217 268
rect 1198 252 1201 258
rect 1210 248 1214 251
rect 1070 132 1073 138
rect 1086 132 1089 148
rect 1110 142 1113 168
rect 1118 132 1121 148
rect 1126 142 1129 218
rect 1158 172 1161 228
rect 1190 192 1193 238
rect 1138 158 1142 161
rect 1150 142 1153 148
rect 838 128 849 131
rect 834 88 838 91
rect 806 62 809 68
rect 846 52 849 128
rect 866 128 870 131
rect 854 92 857 128
rect 878 122 881 128
rect 870 72 873 108
rect 896 103 898 107
rect 902 103 905 107
rect 909 103 912 107
rect 918 72 921 78
rect 914 68 918 71
rect 866 58 870 61
rect 930 58 934 61
rect 878 52 881 58
rect 942 52 945 88
rect 998 72 1001 78
rect 1030 72 1033 78
rect 1018 68 1022 71
rect 974 62 977 68
rect 1038 62 1041 108
rect 1134 92 1137 128
rect 1142 82 1145 138
rect 1114 78 1118 81
rect 1106 68 1110 71
rect 1086 62 1089 68
rect 1010 58 1014 61
rect 1110 52 1113 68
rect 1026 48 1030 51
rect 1058 48 1062 51
rect 862 42 865 48
rect 1126 42 1129 68
rect 1142 62 1145 78
rect 1166 62 1169 188
rect 1190 142 1193 168
rect 1214 162 1217 188
rect 1230 172 1233 228
rect 1238 182 1241 268
rect 1254 192 1257 238
rect 1262 232 1265 258
rect 1246 182 1249 188
rect 1238 172 1241 178
rect 1254 168 1262 171
rect 1226 158 1230 161
rect 1254 151 1257 168
rect 1242 148 1257 151
rect 1262 152 1265 158
rect 1198 142 1201 148
rect 1250 138 1254 141
rect 1174 92 1177 128
rect 1174 72 1177 88
rect 1214 72 1217 118
rect 1230 82 1233 88
rect 1270 62 1273 268
rect 1278 171 1281 268
rect 1298 258 1302 261
rect 1310 252 1313 258
rect 1290 248 1294 251
rect 1318 242 1321 278
rect 1334 272 1337 298
rect 1358 281 1361 368
rect 1350 278 1361 281
rect 1350 252 1353 278
rect 1382 272 1385 338
rect 1358 232 1361 258
rect 1306 218 1310 221
rect 1278 168 1289 171
rect 1278 92 1281 158
rect 1286 152 1289 168
rect 1306 158 1310 161
rect 1318 152 1321 188
rect 1330 178 1334 181
rect 1338 158 1342 161
rect 1306 138 1310 141
rect 1286 132 1289 138
rect 1318 132 1321 138
rect 1326 112 1329 158
rect 1350 152 1353 228
rect 1366 212 1369 268
rect 1374 142 1377 268
rect 1390 262 1393 438
rect 1398 382 1401 468
rect 1406 392 1409 458
rect 1438 452 1441 538
rect 1478 532 1481 538
rect 1462 492 1465 498
rect 1470 481 1473 528
rect 1494 492 1497 648
rect 1502 632 1505 708
rect 1510 692 1513 838
rect 1534 792 1537 958
rect 1542 942 1545 1038
rect 1598 1032 1601 1048
rect 1574 992 1577 1008
rect 1590 992 1593 1028
rect 1630 992 1633 1068
rect 1654 1062 1657 1168
rect 1662 1162 1665 1188
rect 1670 1152 1673 1158
rect 1670 1122 1673 1128
rect 1686 1082 1689 1288
rect 1694 1262 1697 1318
rect 1710 1292 1713 1308
rect 1726 1271 1729 1388
rect 1750 1352 1753 1418
rect 1738 1348 1742 1351
rect 1734 1338 1742 1341
rect 1734 1322 1737 1338
rect 1750 1322 1753 1338
rect 1722 1268 1729 1271
rect 1702 1262 1705 1268
rect 1694 1152 1697 1258
rect 1710 1152 1713 1268
rect 1694 1122 1697 1138
rect 1702 1102 1705 1148
rect 1718 1142 1721 1268
rect 1734 1262 1737 1308
rect 1758 1262 1761 1468
rect 1766 1362 1769 1478
rect 1774 1392 1777 1518
rect 1782 1462 1785 1678
rect 1814 1662 1817 1718
rect 1928 1703 1930 1707
rect 1934 1703 1937 1707
rect 1941 1703 1944 1707
rect 1830 1692 1833 1698
rect 1850 1688 1854 1691
rect 1862 1682 1865 1698
rect 1914 1688 1918 1691
rect 1874 1678 1878 1681
rect 1822 1672 1825 1678
rect 1838 1672 1841 1678
rect 1790 1652 1793 1658
rect 1798 1642 1801 1648
rect 1814 1642 1817 1648
rect 1862 1632 1865 1658
rect 1886 1652 1889 1668
rect 1814 1592 1817 1608
rect 1838 1562 1841 1568
rect 1790 1552 1793 1558
rect 1830 1552 1833 1558
rect 1838 1552 1841 1558
rect 1810 1548 1814 1551
rect 1798 1542 1801 1548
rect 1854 1541 1857 1618
rect 1862 1562 1865 1628
rect 1910 1622 1913 1658
rect 1918 1652 1921 1668
rect 1926 1562 1929 1648
rect 1934 1612 1937 1688
rect 1942 1642 1945 1658
rect 1950 1592 1953 1818
rect 1958 1772 1961 1828
rect 1990 1822 1993 1918
rect 1998 1892 2001 1918
rect 2054 1912 2057 1918
rect 2022 1892 2025 1898
rect 2010 1878 2014 1881
rect 2054 1872 2057 1878
rect 2026 1868 2030 1871
rect 1982 1772 1985 1778
rect 2014 1762 2017 1868
rect 2034 1858 2038 1861
rect 2054 1852 2057 1858
rect 2062 1782 2065 1868
rect 2070 1812 2073 1948
rect 2078 1822 2081 1928
rect 2094 1872 2097 1878
rect 2098 1858 2102 1861
rect 2086 1852 2089 1858
rect 2078 1802 2081 1818
rect 2110 1782 2113 2058
rect 2142 2052 2145 2158
rect 2158 2112 2161 2148
rect 2166 2142 2169 2168
rect 2174 2152 2177 2298
rect 2214 2282 2217 2338
rect 2246 2332 2249 2378
rect 2226 2328 2230 2331
rect 2258 2318 2262 2321
rect 2262 2302 2265 2318
rect 2230 2252 2233 2268
rect 2262 2231 2265 2250
rect 2174 2132 2177 2138
rect 2150 2108 2158 2111
rect 2150 2102 2153 2108
rect 2150 2062 2153 2098
rect 2182 2092 2185 2198
rect 2210 2188 2214 2191
rect 2214 2162 2217 2168
rect 2198 2152 2201 2158
rect 2214 2132 2217 2158
rect 2158 2062 2161 2068
rect 2130 2048 2134 2051
rect 2166 1952 2169 2058
rect 2198 2002 2201 2118
rect 2230 2112 2233 2118
rect 2246 2092 2249 2148
rect 2258 2138 2262 2141
rect 2270 2132 2273 2258
rect 2278 2192 2281 2388
rect 2302 2272 2305 2368
rect 2342 2352 2345 2528
rect 2350 2492 2353 2518
rect 2366 2492 2369 2518
rect 2382 2502 2385 2518
rect 2374 2462 2377 2468
rect 2390 2452 2393 2528
rect 2438 2521 2441 2548
rect 2454 2542 2457 2558
rect 2430 2518 2441 2521
rect 2462 2522 2465 2658
rect 2470 2552 2473 2658
rect 2486 2642 2489 2648
rect 2502 2612 2505 2618
rect 2486 2572 2489 2588
rect 2402 2478 2406 2481
rect 2350 2412 2353 2448
rect 2358 2442 2361 2448
rect 2390 2360 2393 2379
rect 2406 2352 2409 2448
rect 2414 2442 2417 2518
rect 2430 2402 2433 2518
rect 2478 2512 2481 2558
rect 2486 2542 2489 2568
rect 2498 2558 2502 2561
rect 2510 2552 2513 2598
rect 2518 2592 2521 3018
rect 2526 2872 2529 2878
rect 2542 2872 2545 2988
rect 2566 2982 2569 3128
rect 2638 3102 2641 3128
rect 2952 3103 2954 3107
rect 2958 3103 2961 3107
rect 2965 3103 2968 3107
rect 3976 3103 3978 3107
rect 3982 3103 3985 3107
rect 3989 3103 3992 3107
rect 3858 3088 3862 3091
rect 3554 3078 3558 3081
rect 2662 3062 2665 3068
rect 2606 3052 2609 3058
rect 2606 3032 2609 3048
rect 2670 3012 2673 3068
rect 2726 3022 2729 3058
rect 2570 2968 2574 2971
rect 2606 2962 2609 2988
rect 2726 2962 2729 3018
rect 2750 3002 2753 3018
rect 2802 2968 2806 2971
rect 2758 2952 2761 2958
rect 2602 2948 2606 2951
rect 2558 2932 2561 2938
rect 2566 2922 2569 2948
rect 2654 2942 2657 2948
rect 2766 2932 2769 2968
rect 2582 2922 2585 2928
rect 2670 2922 2673 2928
rect 2782 2922 2785 2938
rect 2798 2932 2801 2948
rect 2814 2932 2817 2998
rect 2810 2928 2814 2931
rect 2746 2918 2750 2921
rect 2822 2902 2825 2958
rect 2830 2902 2833 3078
rect 2846 3021 2849 3068
rect 2898 3058 2902 3061
rect 2954 3058 2958 3061
rect 2878 3022 2881 3050
rect 2846 3018 2857 3021
rect 2854 2992 2857 3018
rect 2870 2962 2873 2968
rect 2838 2932 2841 2938
rect 2630 2882 2633 2888
rect 2838 2882 2841 2928
rect 2846 2922 2849 2938
rect 2570 2878 2574 2881
rect 2526 2862 2529 2868
rect 2550 2862 2553 2878
rect 2614 2872 2617 2878
rect 2534 2852 2537 2858
rect 2562 2768 2566 2771
rect 2558 2758 2574 2761
rect 2534 2742 2537 2748
rect 2542 2742 2545 2748
rect 2530 2728 2537 2731
rect 2502 2542 2505 2548
rect 2510 2502 2513 2538
rect 2526 2501 2529 2698
rect 2534 2682 2537 2728
rect 2542 2712 2545 2738
rect 2558 2732 2561 2758
rect 2582 2752 2585 2868
rect 2602 2858 2606 2861
rect 2590 2822 2593 2858
rect 2590 2762 2593 2768
rect 2598 2752 2601 2858
rect 2634 2848 2638 2851
rect 2606 2792 2609 2818
rect 2622 2772 2625 2848
rect 2654 2792 2657 2858
rect 2662 2772 2665 2868
rect 2670 2812 2673 2818
rect 2750 2792 2753 2878
rect 2766 2792 2769 2868
rect 2814 2862 2817 2878
rect 2862 2872 2865 2958
rect 2874 2948 2878 2951
rect 2886 2922 2889 2938
rect 2894 2882 2897 3058
rect 2966 3031 2969 3050
rect 2998 3022 3001 3068
rect 2902 2972 2905 2978
rect 2974 2952 2977 2958
rect 2910 2942 2913 2948
rect 2998 2942 3001 2948
rect 2906 2928 2910 2931
rect 2842 2868 2846 2871
rect 2858 2858 2862 2861
rect 2814 2822 2817 2848
rect 2634 2768 2649 2771
rect 2646 2761 2649 2768
rect 2750 2762 2753 2768
rect 2646 2758 2673 2761
rect 2574 2742 2577 2748
rect 2566 2732 2569 2738
rect 2582 2712 2585 2748
rect 2598 2722 2601 2728
rect 2622 2702 2625 2728
rect 2542 2662 2545 2698
rect 2582 2682 2585 2688
rect 2598 2672 2601 2688
rect 2534 2542 2537 2548
rect 2550 2542 2553 2548
rect 2558 2542 2561 2568
rect 2582 2562 2585 2668
rect 2638 2662 2641 2758
rect 2670 2752 2673 2758
rect 2798 2752 2801 2758
rect 2678 2748 2686 2751
rect 2738 2748 2745 2751
rect 2654 2742 2657 2748
rect 2662 2742 2665 2748
rect 2678 2692 2681 2748
rect 2686 2742 2689 2748
rect 2694 2742 2697 2748
rect 2722 2738 2726 2741
rect 2686 2682 2689 2728
rect 2702 2712 2705 2738
rect 2722 2728 2726 2731
rect 2682 2678 2686 2681
rect 2694 2672 2697 2698
rect 2710 2672 2713 2718
rect 2734 2682 2737 2688
rect 2742 2672 2745 2748
rect 2826 2748 2830 2751
rect 2750 2742 2753 2748
rect 2782 2742 2785 2748
rect 2802 2738 2806 2741
rect 2758 2732 2761 2738
rect 2750 2722 2753 2728
rect 2774 2692 2777 2728
rect 2790 2722 2793 2738
rect 2814 2682 2817 2748
rect 2830 2702 2833 2738
rect 2838 2712 2841 2738
rect 2846 2722 2849 2728
rect 2722 2668 2726 2671
rect 2754 2668 2758 2671
rect 2722 2658 2734 2661
rect 2670 2652 2673 2658
rect 2630 2631 2633 2650
rect 2638 2592 2641 2648
rect 2670 2592 2673 2638
rect 2586 2558 2590 2561
rect 2654 2552 2657 2558
rect 2542 2522 2545 2538
rect 2570 2518 2574 2521
rect 2598 2502 2601 2548
rect 2606 2542 2609 2548
rect 2618 2528 2622 2531
rect 2650 2528 2654 2531
rect 2670 2522 2673 2548
rect 2686 2542 2689 2648
rect 2702 2642 2705 2658
rect 2742 2652 2745 2668
rect 2766 2662 2769 2668
rect 2750 2652 2753 2658
rect 2718 2622 2721 2648
rect 2718 2602 2721 2618
rect 2790 2582 2793 2658
rect 2802 2648 2806 2651
rect 2818 2618 2822 2621
rect 2822 2560 2825 2579
rect 2686 2511 2689 2538
rect 2698 2518 2702 2521
rect 2686 2508 2697 2511
rect 2526 2498 2537 2501
rect 2486 2472 2489 2478
rect 2502 2472 2505 2488
rect 2534 2462 2537 2498
rect 2578 2478 2582 2481
rect 2598 2478 2606 2481
rect 2582 2472 2585 2478
rect 2598 2472 2601 2478
rect 2614 2472 2617 2508
rect 2626 2488 2630 2491
rect 2606 2462 2609 2468
rect 2630 2461 2633 2478
rect 2646 2462 2649 2468
rect 2630 2458 2638 2461
rect 2446 2452 2449 2458
rect 2590 2452 2593 2458
rect 2618 2448 2622 2451
rect 2440 2403 2442 2407
rect 2446 2403 2449 2407
rect 2453 2403 2456 2407
rect 2486 2392 2489 2448
rect 2358 2342 2361 2348
rect 2342 2332 2345 2338
rect 2342 2311 2345 2318
rect 2326 2308 2345 2311
rect 2326 2292 2329 2308
rect 2334 2272 2337 2278
rect 2302 2202 2305 2268
rect 2350 2262 2353 2268
rect 2366 2262 2369 2298
rect 2390 2282 2393 2338
rect 2402 2278 2406 2281
rect 2414 2272 2417 2378
rect 2502 2362 2505 2438
rect 2550 2422 2553 2448
rect 2566 2372 2569 2418
rect 2474 2358 2478 2361
rect 2518 2352 2521 2358
rect 2542 2352 2545 2368
rect 2566 2362 2569 2368
rect 2466 2348 2470 2351
rect 2454 2342 2457 2348
rect 2478 2342 2481 2348
rect 2518 2342 2521 2348
rect 2526 2342 2529 2348
rect 2574 2342 2577 2418
rect 2654 2382 2657 2468
rect 2662 2462 2665 2508
rect 2694 2492 2697 2508
rect 2710 2492 2713 2498
rect 2718 2472 2721 2558
rect 2774 2532 2777 2548
rect 2790 2532 2793 2538
rect 2734 2472 2737 2478
rect 2774 2472 2777 2498
rect 2830 2492 2833 2698
rect 2838 2622 2841 2708
rect 2862 2702 2865 2758
rect 2878 2742 2881 2748
rect 2886 2742 2889 2748
rect 2902 2682 2905 2898
rect 2942 2892 2945 2918
rect 2952 2903 2954 2907
rect 2958 2903 2961 2907
rect 2965 2903 2968 2907
rect 2934 2832 2937 2878
rect 2950 2862 2953 2868
rect 2982 2862 2985 2878
rect 3002 2818 3006 2821
rect 2918 2792 2921 2818
rect 3014 2802 3017 3078
rect 3054 3042 3057 3078
rect 3122 3058 3126 3061
rect 3054 2992 3057 3038
rect 3086 2992 3089 3058
rect 3098 3028 3102 3031
rect 3070 2942 3073 2948
rect 3102 2922 3105 2948
rect 3118 2932 3121 2948
rect 3054 2902 3057 2918
rect 3110 2902 3113 2918
rect 3078 2882 3081 2898
rect 3126 2892 3129 2938
rect 3094 2872 3097 2878
rect 3134 2862 3137 3058
rect 3142 3022 3145 3050
rect 3174 3021 3177 3068
rect 3190 3042 3193 3078
rect 3298 3058 3302 3061
rect 3166 3018 3177 3021
rect 3166 2992 3169 3018
rect 3198 2992 3201 3018
rect 3142 2952 3145 2958
rect 3162 2948 3166 2951
rect 3126 2831 3129 2850
rect 3134 2802 3137 2858
rect 3142 2852 3145 2948
rect 3166 2872 3169 2938
rect 2918 2772 2921 2788
rect 2958 2732 2961 2748
rect 2998 2732 3001 2798
rect 3014 2742 3017 2768
rect 3046 2760 3049 2779
rect 3062 2752 3065 2798
rect 3098 2768 3102 2771
rect 3126 2752 3129 2758
rect 3134 2752 3137 2798
rect 3166 2782 3169 2868
rect 3174 2802 3177 2938
rect 3182 2892 3185 2958
rect 3194 2948 3198 2951
rect 3206 2942 3209 2968
rect 3230 2952 3233 3058
rect 3302 3022 3305 3048
rect 3270 2992 3273 3018
rect 3246 2960 3249 2979
rect 3190 2862 3193 2898
rect 3206 2892 3209 2928
rect 3198 2862 3201 2868
rect 3214 2852 3217 2868
rect 3222 2862 3225 2948
rect 3278 2932 3281 2938
rect 3294 2932 3297 2958
rect 3278 2882 3281 2918
rect 3334 2902 3337 2948
rect 3350 2902 3353 3068
rect 3366 3052 3369 3078
rect 3494 3042 3497 3058
rect 3502 3052 3505 3078
rect 3518 3062 3521 3068
rect 3570 3058 3574 3061
rect 3526 3042 3529 3058
rect 3550 3052 3553 3058
rect 3590 3052 3593 3078
rect 3614 3072 3617 3088
rect 3646 3072 3649 3088
rect 4094 3082 4097 3088
rect 4262 3082 4265 3088
rect 3674 3078 3678 3081
rect 3850 3078 3854 3081
rect 4290 3078 4294 3081
rect 3618 3058 3622 3061
rect 3618 3048 3622 3051
rect 3450 3018 3454 3021
rect 3472 3003 3474 3007
rect 3478 3003 3481 3007
rect 3485 3003 3488 3007
rect 3438 2962 3441 2978
rect 3446 2962 3449 2968
rect 3494 2962 3497 3018
rect 3502 3012 3505 3038
rect 3518 3012 3521 3038
rect 3566 3032 3569 3038
rect 3558 2992 3561 3028
rect 3482 2958 3486 2961
rect 3422 2952 3425 2958
rect 3430 2952 3433 2958
rect 3406 2942 3409 2948
rect 3438 2942 3441 2948
rect 3386 2928 3390 2931
rect 3418 2928 3422 2931
rect 3370 2918 3374 2921
rect 3374 2912 3377 2918
rect 3230 2852 3233 2878
rect 3278 2872 3281 2878
rect 3270 2862 3273 2868
rect 3318 2862 3321 2898
rect 3350 2862 3353 2868
rect 3242 2858 3246 2861
rect 3186 2848 3190 2851
rect 3254 2832 3257 2858
rect 3262 2852 3265 2858
rect 3302 2822 3305 2848
rect 3366 2792 3369 2878
rect 3406 2812 3409 2928
rect 3478 2892 3481 2948
rect 3558 2942 3561 2988
rect 3566 2972 3569 2978
rect 3494 2892 3497 2928
rect 3502 2922 3505 2938
rect 3534 2902 3537 2918
rect 3550 2912 3553 2938
rect 3502 2892 3505 2898
rect 3518 2882 3521 2888
rect 3450 2818 3454 2821
rect 3446 2792 3449 2808
rect 3190 2760 3193 2779
rect 3322 2778 3326 2781
rect 3434 2768 3438 2771
rect 3450 2768 3454 2771
rect 3462 2771 3465 2868
rect 3502 2862 3505 2878
rect 3526 2871 3529 2888
rect 3558 2882 3561 2888
rect 3546 2878 3550 2881
rect 3514 2868 3529 2871
rect 3566 2871 3569 2948
rect 3574 2892 3577 3018
rect 3582 2982 3585 3048
rect 3654 3042 3657 3068
rect 3670 3062 3673 3068
rect 3686 3052 3689 3068
rect 3694 3062 3697 3068
rect 3702 3062 3705 3068
rect 3670 3042 3673 3048
rect 3702 3042 3705 3058
rect 3718 3042 3721 3078
rect 3750 3072 3753 3078
rect 3766 3072 3769 3078
rect 3742 3062 3745 3068
rect 3790 3062 3793 3068
rect 3822 3062 3825 3068
rect 3758 3052 3761 3058
rect 3766 3052 3769 3058
rect 3794 3048 3798 3051
rect 3606 3022 3609 3028
rect 3654 3022 3657 3038
rect 3638 2962 3641 3018
rect 3670 2992 3673 3028
rect 3582 2892 3585 2958
rect 3614 2952 3617 2958
rect 3590 2932 3593 2948
rect 3622 2942 3625 2958
rect 3670 2952 3673 2988
rect 3694 2961 3697 2978
rect 3694 2958 3702 2961
rect 3658 2948 3662 2951
rect 3678 2932 3681 2938
rect 3694 2932 3697 2958
rect 3710 2952 3713 2998
rect 3718 2992 3721 3008
rect 3718 2972 3721 2988
rect 3742 2972 3745 3018
rect 3758 2992 3761 3048
rect 3774 3042 3777 3048
rect 3766 2992 3769 3038
rect 3766 2982 3769 2988
rect 3754 2968 3758 2971
rect 3782 2962 3785 3048
rect 3814 3012 3817 3048
rect 3822 3042 3825 3058
rect 3830 3042 3833 3048
rect 3822 2992 3825 3018
rect 3830 2992 3833 3038
rect 3802 2968 3806 2971
rect 3734 2932 3737 2958
rect 3690 2928 3694 2931
rect 3590 2881 3593 2928
rect 3638 2922 3641 2928
rect 3630 2902 3633 2918
rect 3582 2878 3593 2881
rect 3566 2868 3574 2871
rect 3550 2862 3553 2868
rect 3574 2862 3577 2868
rect 3490 2858 3494 2861
rect 3494 2812 3497 2848
rect 3472 2803 3474 2807
rect 3478 2803 3481 2807
rect 3485 2803 3488 2807
rect 3506 2788 3510 2791
rect 3462 2768 3470 2771
rect 3470 2762 3473 2768
rect 3518 2752 3521 2848
rect 3542 2842 3545 2858
rect 3550 2802 3553 2858
rect 3566 2792 3569 2858
rect 3574 2842 3577 2858
rect 3582 2762 3585 2878
rect 3598 2872 3601 2878
rect 3618 2858 3622 2861
rect 3590 2822 3593 2848
rect 3078 2748 3086 2751
rect 3170 2748 3174 2751
rect 3394 2748 3398 2751
rect 3442 2748 3446 2751
rect 2998 2722 3001 2728
rect 2914 2718 2918 2721
rect 2952 2703 2954 2707
rect 2958 2703 2961 2707
rect 2965 2703 2968 2707
rect 3030 2682 3033 2688
rect 2842 2548 2846 2551
rect 2814 2472 2817 2488
rect 2698 2468 2702 2471
rect 2802 2468 2806 2471
rect 2678 2462 2681 2468
rect 2686 2432 2689 2468
rect 2718 2392 2721 2468
rect 2730 2458 2734 2461
rect 2742 2452 2745 2468
rect 2750 2462 2753 2468
rect 2854 2462 2857 2608
rect 2754 2448 2758 2451
rect 2750 2392 2753 2428
rect 2586 2368 2590 2371
rect 2634 2368 2638 2371
rect 2606 2362 2609 2368
rect 2654 2362 2657 2368
rect 2662 2362 2665 2368
rect 2678 2352 2681 2388
rect 2766 2372 2769 2428
rect 2774 2392 2777 2458
rect 2782 2452 2785 2458
rect 2790 2362 2793 2408
rect 2806 2372 2809 2378
rect 2774 2352 2777 2358
rect 2738 2348 2742 2351
rect 2590 2342 2593 2348
rect 2638 2342 2641 2348
rect 2790 2342 2793 2348
rect 2798 2342 2801 2358
rect 2814 2352 2817 2458
rect 2846 2422 2849 2458
rect 2822 2352 2825 2388
rect 2838 2362 2841 2398
rect 2854 2392 2857 2448
rect 2862 2362 2865 2528
rect 2902 2512 2905 2678
rect 3014 2672 3017 2678
rect 3002 2668 3006 2671
rect 3034 2668 3038 2671
rect 2918 2612 2921 2668
rect 2950 2662 2953 2668
rect 3022 2662 3025 2668
rect 3046 2662 3049 2698
rect 3066 2668 3070 2671
rect 3078 2662 3081 2748
rect 3110 2742 3113 2748
rect 3130 2738 3134 2741
rect 3086 2692 3089 2738
rect 3094 2692 3097 2728
rect 3118 2712 3121 2738
rect 3142 2692 3145 2748
rect 3222 2742 3225 2748
rect 3102 2672 3105 2688
rect 3094 2662 3097 2668
rect 3110 2662 3113 2668
rect 3066 2658 3070 2661
rect 3082 2658 3089 2661
rect 3122 2658 3126 2661
rect 2966 2622 2969 2648
rect 3062 2642 3065 2648
rect 3086 2642 3089 2658
rect 3134 2652 3137 2668
rect 3150 2652 3153 2738
rect 3238 2732 3241 2738
rect 3254 2692 3257 2708
rect 3190 2682 3193 2688
rect 3262 2682 3265 2688
rect 3278 2682 3281 2748
rect 3382 2742 3385 2748
rect 3362 2718 3366 2721
rect 3382 2712 3385 2738
rect 3398 2722 3401 2738
rect 3406 2732 3409 2738
rect 3418 2728 3422 2731
rect 3462 2722 3465 2748
rect 3494 2732 3497 2738
rect 3502 2712 3505 2748
rect 3166 2672 3169 2678
rect 3286 2672 3289 2688
rect 3430 2682 3433 2688
rect 3162 2658 3166 2661
rect 3110 2642 3113 2648
rect 3014 2562 3017 2588
rect 2910 2542 2913 2548
rect 2966 2542 2969 2548
rect 3006 2542 3009 2548
rect 2910 2472 2913 2528
rect 2950 2522 2953 2528
rect 2926 2472 2929 2478
rect 2874 2458 2878 2461
rect 2894 2442 2897 2468
rect 2906 2458 2910 2461
rect 2870 2382 2873 2418
rect 2902 2362 2905 2458
rect 2918 2452 2921 2458
rect 2934 2392 2937 2508
rect 2952 2503 2954 2507
rect 2958 2503 2961 2507
rect 2965 2503 2968 2507
rect 2958 2462 2961 2488
rect 2982 2462 2985 2468
rect 3006 2462 3009 2468
rect 3030 2462 3033 2558
rect 3054 2542 3057 2578
rect 3062 2531 3065 2638
rect 3086 2592 3089 2638
rect 3142 2632 3145 2648
rect 3174 2642 3177 2658
rect 3110 2592 3113 2608
rect 3086 2582 3089 2588
rect 3146 2568 3150 2571
rect 3054 2528 3065 2531
rect 3146 2548 3150 2551
rect 3038 2462 3041 2468
rect 2950 2422 2953 2458
rect 2998 2422 3001 2458
rect 2974 2402 2977 2418
rect 3022 2382 3025 2418
rect 2874 2358 2878 2361
rect 2578 2338 2582 2341
rect 2682 2338 2686 2341
rect 2754 2338 2758 2341
rect 2446 2322 2449 2338
rect 2454 2282 2457 2288
rect 2398 2268 2414 2271
rect 2450 2268 2454 2271
rect 2390 2262 2393 2268
rect 2314 2258 2318 2261
rect 2338 2258 2342 2261
rect 2382 2242 2385 2248
rect 2278 2182 2281 2188
rect 2318 2162 2321 2168
rect 2326 2152 2329 2178
rect 2366 2162 2369 2188
rect 2298 2148 2302 2151
rect 2350 2142 2353 2158
rect 2290 2138 2294 2141
rect 2330 2138 2334 2141
rect 2318 2102 2321 2118
rect 2286 2082 2289 2098
rect 2302 2062 2305 2068
rect 2334 2062 2337 2128
rect 2350 2062 2353 2118
rect 2358 2112 2361 2148
rect 2382 2142 2385 2238
rect 2398 2201 2401 2268
rect 2422 2262 2425 2268
rect 2470 2262 2473 2308
rect 2410 2258 2422 2261
rect 2440 2203 2442 2207
rect 2446 2203 2449 2207
rect 2453 2203 2456 2207
rect 2394 2198 2401 2201
rect 2390 2142 2393 2198
rect 2478 2182 2481 2338
rect 2534 2332 2537 2338
rect 2562 2328 2566 2331
rect 2550 2282 2553 2308
rect 2494 2272 2497 2278
rect 2554 2268 2558 2271
rect 2506 2248 2510 2251
rect 2486 2242 2489 2248
rect 2418 2158 2422 2161
rect 2490 2148 2494 2151
rect 2382 2132 2385 2138
rect 2398 2102 2401 2148
rect 2430 2132 2433 2138
rect 2382 2092 2385 2098
rect 2406 2092 2409 2108
rect 2414 2082 2417 2118
rect 2438 2112 2441 2148
rect 2446 2142 2449 2148
rect 2502 2142 2505 2198
rect 2526 2182 2529 2268
rect 2574 2262 2577 2318
rect 2614 2302 2617 2328
rect 2586 2268 2590 2271
rect 2606 2262 2609 2268
rect 2630 2262 2633 2338
rect 2558 2258 2566 2261
rect 2578 2258 2582 2261
rect 2594 2258 2598 2261
rect 2558 2251 2561 2258
rect 2554 2248 2561 2251
rect 2570 2248 2577 2251
rect 2574 2232 2577 2248
rect 2386 2078 2390 2081
rect 2454 2072 2457 2138
rect 2534 2132 2537 2138
rect 2466 2128 2470 2131
rect 2506 2128 2513 2131
rect 2538 2128 2542 2131
rect 2470 2072 2473 2098
rect 2502 2072 2505 2078
rect 2510 2072 2513 2128
rect 2526 2092 2529 2098
rect 2550 2082 2553 2178
rect 2566 2162 2569 2228
rect 2574 2192 2577 2228
rect 2590 2152 2593 2258
rect 2638 2252 2641 2338
rect 2694 2332 2697 2338
rect 2766 2332 2769 2338
rect 2706 2328 2710 2331
rect 2822 2322 2825 2348
rect 2838 2342 2841 2348
rect 2846 2342 2849 2348
rect 2854 2332 2857 2348
rect 2878 2342 2881 2348
rect 2886 2342 2889 2348
rect 2910 2342 2913 2368
rect 3002 2358 3006 2361
rect 2898 2338 2902 2341
rect 2662 2282 2665 2318
rect 2750 2312 2753 2318
rect 2830 2292 2833 2318
rect 2926 2282 2929 2358
rect 2998 2352 3001 2358
rect 3014 2352 3017 2368
rect 2934 2342 2937 2348
rect 2990 2342 2993 2348
rect 3022 2342 3025 2348
rect 2970 2328 2974 2331
rect 2952 2303 2954 2307
rect 2958 2303 2961 2307
rect 2965 2303 2968 2307
rect 2734 2272 2737 2278
rect 2942 2272 2945 2278
rect 2650 2218 2654 2221
rect 2622 2212 2625 2218
rect 2562 2148 2566 2151
rect 2590 2142 2593 2148
rect 2578 2138 2582 2141
rect 2558 2122 2561 2128
rect 2598 2112 2601 2148
rect 2638 2142 2641 2218
rect 2678 2152 2681 2158
rect 2654 2142 2657 2148
rect 2686 2142 2689 2148
rect 2694 2142 2697 2198
rect 2722 2188 2726 2191
rect 2726 2182 2729 2188
rect 2630 2132 2633 2138
rect 2682 2118 2686 2121
rect 2646 2102 2649 2118
rect 2622 2082 2625 2088
rect 2638 2072 2641 2098
rect 2426 2068 2430 2071
rect 2370 2058 2374 2061
rect 2206 2012 2209 2018
rect 2334 2011 2337 2058
rect 2350 2022 2353 2048
rect 2326 2008 2337 2011
rect 2230 1962 2233 1988
rect 2326 1952 2329 2008
rect 2366 1952 2369 2058
rect 2398 2012 2401 2068
rect 2438 2062 2441 2068
rect 2418 2058 2422 2061
rect 2478 2032 2481 2058
rect 2494 2052 2497 2058
rect 2440 2003 2442 2007
rect 2446 2003 2449 2007
rect 2453 2003 2456 2007
rect 2430 1962 2433 1988
rect 2510 1962 2513 2058
rect 2582 2052 2585 2058
rect 2530 2048 2534 2051
rect 2538 2028 2542 2031
rect 2478 1952 2481 1958
rect 2274 1948 2278 1951
rect 2498 1948 2502 1951
rect 2514 1948 2518 1951
rect 2126 1911 2129 1948
rect 2230 1942 2233 1948
rect 2326 1942 2329 1948
rect 2382 1942 2385 1948
rect 2166 1932 2169 1938
rect 2182 1922 2185 1938
rect 2366 1932 2369 1938
rect 2250 1928 2254 1931
rect 2118 1908 2129 1911
rect 2118 1892 2121 1908
rect 2126 1862 2129 1898
rect 2134 1862 2137 1908
rect 2182 1862 2185 1888
rect 2222 1882 2225 1928
rect 2278 1922 2281 1928
rect 2262 1912 2265 1918
rect 2230 1882 2233 1888
rect 2218 1878 2222 1881
rect 2146 1858 2150 1861
rect 2162 1848 2166 1851
rect 2174 1802 2177 1858
rect 2198 1842 2201 1868
rect 2246 1862 2249 1868
rect 2258 1866 2262 1869
rect 2070 1762 2073 1768
rect 2082 1758 2086 1761
rect 1998 1742 2001 1748
rect 1986 1738 1990 1741
rect 2006 1738 2022 1741
rect 1958 1692 1961 1698
rect 1958 1622 1961 1628
rect 1966 1611 1969 1728
rect 1990 1692 1993 1728
rect 1998 1702 2001 1738
rect 2006 1712 2009 1738
rect 2030 1732 2033 1748
rect 2046 1732 2049 1748
rect 2054 1742 2057 1758
rect 2110 1752 2113 1778
rect 2158 1762 2161 1768
rect 2182 1762 2185 1778
rect 2190 1771 2193 1818
rect 2190 1768 2201 1771
rect 2146 1758 2150 1761
rect 2190 1752 2193 1758
rect 2062 1742 2065 1748
rect 2070 1742 2073 1748
rect 2018 1728 2022 1731
rect 1974 1632 1977 1668
rect 2014 1662 2017 1698
rect 2022 1682 2025 1708
rect 2030 1672 2033 1718
rect 2038 1672 2041 1708
rect 2054 1672 2057 1698
rect 2062 1662 2065 1668
rect 2070 1662 2073 1738
rect 2086 1732 2089 1748
rect 2198 1742 2201 1768
rect 2206 1752 2209 1858
rect 2218 1848 2222 1851
rect 2238 1851 2241 1858
rect 2238 1848 2254 1851
rect 2278 1812 2281 1918
rect 2430 1912 2433 1948
rect 2486 1942 2489 1948
rect 2506 1938 2513 1941
rect 2462 1922 2465 1938
rect 2294 1872 2297 1908
rect 2290 1858 2294 1861
rect 2302 1852 2305 1888
rect 2358 1882 2361 1908
rect 2378 1888 2382 1891
rect 2398 1882 2401 1888
rect 2334 1862 2337 1868
rect 2314 1858 2318 1861
rect 2270 1762 2273 1768
rect 2218 1758 2222 1761
rect 2242 1758 2246 1761
rect 2310 1752 2313 1848
rect 2326 1822 2329 1858
rect 2342 1852 2345 1858
rect 2358 1772 2361 1878
rect 2366 1862 2369 1868
rect 2382 1852 2385 1858
rect 2390 1822 2393 1878
rect 2406 1862 2409 1868
rect 2406 1842 2409 1848
rect 2414 1752 2417 1908
rect 2430 1872 2433 1878
rect 2438 1862 2441 1898
rect 2454 1872 2457 1918
rect 2462 1892 2465 1918
rect 2502 1872 2505 1908
rect 2510 1872 2513 1938
rect 2534 1932 2537 1938
rect 2542 1921 2545 1958
rect 2534 1918 2545 1921
rect 2502 1862 2505 1868
rect 2474 1858 2478 1861
rect 2534 1842 2537 1918
rect 2550 1862 2553 2048
rect 2670 2031 2673 2050
rect 2558 1952 2561 1968
rect 2566 1922 2569 1938
rect 2574 1932 2577 2028
rect 2614 1992 2617 2008
rect 2646 1992 2649 2008
rect 2666 1988 2670 1991
rect 2582 1972 2585 1978
rect 2590 1952 2593 1958
rect 2622 1952 2625 1968
rect 2634 1958 2638 1961
rect 2598 1942 2601 1948
rect 2658 1938 2662 1941
rect 2654 1902 2657 1938
rect 2590 1882 2593 1888
rect 2678 1882 2681 1888
rect 2606 1872 2609 1878
rect 2678 1862 2681 1868
rect 2546 1858 2550 1861
rect 2506 1818 2510 1821
rect 2440 1803 2442 1807
rect 2446 1803 2449 1807
rect 2453 1803 2456 1807
rect 2422 1762 2425 1788
rect 2478 1762 2481 1768
rect 2462 1752 2465 1758
rect 2162 1738 2166 1741
rect 2186 1738 2190 1741
rect 2218 1738 2222 1741
rect 2098 1728 2102 1731
rect 2118 1692 2121 1728
rect 2106 1688 2110 1691
rect 2126 1682 2129 1718
rect 2134 1712 2137 1728
rect 2142 1702 2145 1738
rect 2230 1732 2233 1748
rect 2250 1738 2254 1741
rect 2274 1718 2278 1721
rect 2174 1681 2177 1718
rect 2246 1702 2249 1718
rect 2278 1712 2281 1718
rect 2166 1678 2177 1681
rect 2262 1682 2265 1688
rect 2086 1662 2089 1678
rect 2130 1668 2134 1671
rect 2154 1668 2158 1671
rect 2110 1662 2113 1668
rect 2026 1658 2030 1661
rect 1998 1632 2001 1648
rect 2070 1642 2073 1648
rect 2058 1618 2062 1621
rect 1958 1608 1969 1611
rect 2094 1612 2097 1648
rect 1862 1552 1865 1558
rect 1950 1552 1953 1558
rect 1898 1548 1902 1551
rect 1870 1542 1873 1548
rect 1854 1538 1862 1541
rect 1898 1538 1902 1541
rect 1806 1472 1809 1538
rect 1838 1482 1841 1518
rect 1846 1482 1849 1508
rect 1870 1491 1873 1538
rect 1910 1531 1913 1548
rect 1946 1538 1950 1541
rect 1902 1528 1913 1531
rect 1862 1488 1873 1491
rect 1822 1472 1825 1478
rect 1830 1472 1833 1478
rect 1814 1462 1817 1468
rect 1826 1458 1830 1461
rect 1798 1452 1801 1458
rect 1770 1348 1774 1351
rect 1818 1348 1822 1351
rect 1778 1318 1782 1321
rect 1790 1302 1793 1348
rect 1806 1322 1809 1328
rect 1814 1302 1817 1338
rect 1830 1312 1833 1448
rect 1854 1402 1857 1458
rect 1846 1362 1849 1388
rect 1838 1332 1841 1358
rect 1854 1352 1857 1398
rect 1862 1362 1865 1488
rect 1870 1452 1873 1478
rect 1878 1392 1881 1468
rect 1882 1358 1886 1361
rect 1894 1352 1897 1518
rect 1902 1492 1905 1528
rect 1958 1522 1961 1608
rect 2018 1588 2022 1591
rect 1982 1562 1985 1568
rect 1966 1552 1969 1558
rect 1998 1552 2001 1558
rect 1928 1503 1930 1507
rect 1934 1503 1937 1507
rect 1941 1503 1944 1507
rect 1974 1492 1977 1538
rect 2006 1532 2009 1588
rect 2022 1542 2025 1548
rect 1930 1478 1934 1481
rect 2030 1472 2033 1558
rect 2054 1552 2057 1588
rect 2070 1561 2073 1568
rect 2062 1558 2073 1561
rect 2062 1552 2065 1558
rect 2042 1518 2046 1521
rect 2070 1512 2073 1548
rect 2086 1532 2089 1598
rect 2118 1572 2121 1648
rect 2142 1642 2145 1668
rect 2166 1661 2169 1678
rect 2154 1658 2169 1661
rect 2174 1652 2177 1668
rect 2278 1642 2281 1668
rect 2318 1662 2321 1748
rect 2358 1732 2361 1738
rect 2374 1732 2377 1738
rect 2478 1712 2481 1748
rect 2166 1592 2169 1638
rect 2154 1558 2158 1561
rect 2122 1548 2126 1551
rect 2122 1538 2126 1541
rect 2078 1528 2086 1531
rect 1902 1462 1905 1468
rect 1998 1462 2001 1468
rect 2038 1462 2041 1498
rect 1914 1458 1918 1461
rect 1970 1458 1974 1461
rect 2018 1458 2022 1461
rect 1902 1382 1905 1388
rect 1874 1348 1878 1351
rect 1898 1348 1902 1351
rect 1846 1332 1849 1348
rect 1886 1322 1889 1338
rect 1766 1272 1769 1278
rect 1742 1192 1745 1218
rect 1734 1162 1737 1168
rect 1726 1132 1729 1158
rect 1742 1132 1745 1188
rect 1758 1171 1761 1258
rect 1754 1168 1761 1171
rect 1766 1161 1769 1218
rect 1774 1202 1777 1278
rect 1782 1262 1785 1268
rect 1814 1262 1817 1288
rect 1822 1262 1825 1268
rect 1794 1258 1798 1261
rect 1834 1258 1838 1261
rect 1854 1261 1857 1318
rect 1854 1258 1862 1261
rect 1798 1192 1801 1258
rect 1850 1228 1854 1231
rect 1758 1158 1769 1161
rect 1758 1152 1761 1158
rect 1814 1152 1817 1188
rect 1878 1182 1881 1278
rect 1886 1261 1889 1308
rect 1894 1302 1897 1338
rect 1902 1272 1905 1338
rect 1886 1258 1894 1261
rect 1910 1252 1913 1258
rect 1910 1192 1913 1218
rect 1918 1192 1921 1398
rect 1958 1372 1961 1458
rect 1990 1442 1993 1458
rect 2006 1431 2009 1448
rect 2022 1442 2025 1448
rect 1998 1428 2009 1431
rect 1962 1358 1969 1361
rect 1926 1342 1929 1358
rect 1966 1352 1969 1358
rect 1926 1332 1929 1338
rect 1928 1303 1930 1307
rect 1934 1303 1937 1307
rect 1941 1303 1944 1307
rect 1950 1291 1953 1328
rect 1946 1288 1953 1291
rect 1958 1272 1961 1348
rect 1934 1252 1937 1268
rect 1946 1258 1950 1261
rect 1826 1148 1830 1151
rect 1722 1128 1726 1131
rect 1750 1122 1753 1128
rect 1758 1111 1761 1148
rect 1790 1142 1793 1148
rect 1822 1132 1825 1138
rect 1830 1132 1833 1148
rect 1750 1108 1761 1111
rect 1638 1042 1641 1058
rect 1650 1048 1654 1051
rect 1574 952 1577 978
rect 1562 948 1569 951
rect 1542 892 1545 928
rect 1542 872 1545 878
rect 1550 872 1553 908
rect 1542 862 1545 868
rect 1558 852 1561 898
rect 1566 841 1569 948
rect 1582 942 1585 948
rect 1602 938 1606 941
rect 1582 892 1585 908
rect 1582 872 1585 888
rect 1598 871 1601 928
rect 1614 922 1617 948
rect 1638 942 1641 958
rect 1642 928 1646 931
rect 1594 868 1601 871
rect 1574 862 1577 868
rect 1558 838 1569 841
rect 1558 792 1561 838
rect 1574 772 1577 818
rect 1582 792 1585 838
rect 1590 792 1593 868
rect 1614 852 1617 898
rect 1662 892 1665 1058
rect 1670 962 1673 1058
rect 1686 1052 1689 1068
rect 1694 1002 1697 1068
rect 1702 1062 1705 1098
rect 1734 1092 1737 1098
rect 1710 1072 1713 1078
rect 1750 1062 1753 1108
rect 1694 952 1697 988
rect 1718 982 1721 1048
rect 1722 958 1726 961
rect 1706 948 1710 951
rect 1646 872 1649 878
rect 1638 862 1641 868
rect 1598 832 1601 838
rect 1638 802 1641 818
rect 1618 778 1622 781
rect 1522 758 1526 761
rect 1546 758 1550 761
rect 1518 722 1521 748
rect 1526 732 1529 738
rect 1526 692 1529 718
rect 1558 691 1561 768
rect 1598 762 1601 768
rect 1626 748 1630 751
rect 1566 702 1569 728
rect 1574 722 1577 738
rect 1550 688 1561 691
rect 1550 672 1553 688
rect 1562 678 1566 681
rect 1518 662 1521 668
rect 1510 572 1513 648
rect 1526 642 1529 658
rect 1518 592 1521 628
rect 1582 592 1585 748
rect 1642 738 1646 741
rect 1630 732 1633 738
rect 1606 712 1609 728
rect 1622 692 1625 728
rect 1638 712 1641 718
rect 1646 712 1649 721
rect 1654 712 1657 878
rect 1670 862 1673 948
rect 1742 932 1745 938
rect 1666 858 1670 861
rect 1662 752 1665 838
rect 1670 792 1673 828
rect 1678 812 1681 918
rect 1702 882 1705 888
rect 1710 872 1713 928
rect 1718 902 1721 928
rect 1726 882 1729 888
rect 1686 862 1689 868
rect 1726 862 1729 878
rect 1734 872 1737 878
rect 1706 858 1710 861
rect 1686 762 1689 768
rect 1670 742 1673 748
rect 1694 742 1697 858
rect 1702 842 1705 848
rect 1702 792 1705 798
rect 1734 792 1737 808
rect 1722 758 1726 761
rect 1730 748 1734 751
rect 1702 742 1705 748
rect 1662 722 1665 738
rect 1646 672 1649 708
rect 1654 682 1657 698
rect 1686 692 1689 738
rect 1726 722 1729 738
rect 1710 678 1737 681
rect 1606 662 1609 668
rect 1614 662 1617 668
rect 1678 662 1681 668
rect 1702 662 1705 678
rect 1710 672 1713 678
rect 1734 672 1737 678
rect 1590 642 1593 648
rect 1502 562 1505 568
rect 1534 562 1537 568
rect 1590 552 1593 608
rect 1614 552 1617 558
rect 1622 552 1625 658
rect 1670 652 1673 658
rect 1630 562 1633 568
rect 1638 552 1641 618
rect 1646 592 1649 608
rect 1506 548 1510 551
rect 1538 548 1542 551
rect 1562 548 1566 551
rect 1510 512 1513 538
rect 1554 528 1558 531
rect 1518 492 1521 528
rect 1566 521 1569 538
rect 1558 518 1569 521
rect 1462 478 1473 481
rect 1482 478 1486 481
rect 1454 472 1457 478
rect 1462 462 1465 478
rect 1474 468 1478 471
rect 1450 458 1454 461
rect 1482 458 1486 461
rect 1416 403 1418 407
rect 1422 403 1425 407
rect 1429 403 1432 407
rect 1454 372 1457 458
rect 1474 358 1478 361
rect 1422 352 1425 358
rect 1486 352 1489 398
rect 1398 272 1401 348
rect 1430 262 1433 348
rect 1442 268 1446 271
rect 1410 258 1414 261
rect 1382 252 1385 258
rect 1422 222 1425 248
rect 1382 152 1385 218
rect 1398 202 1401 218
rect 1416 203 1418 207
rect 1422 203 1425 207
rect 1429 203 1432 207
rect 1358 102 1361 138
rect 1370 128 1374 131
rect 1382 122 1385 138
rect 1390 92 1393 158
rect 1398 152 1401 168
rect 1414 152 1417 158
rect 1438 152 1441 228
rect 1446 202 1449 238
rect 1454 232 1457 348
rect 1494 342 1497 468
rect 1510 462 1513 478
rect 1526 472 1529 478
rect 1534 472 1537 478
rect 1506 368 1510 371
rect 1510 352 1513 358
rect 1474 338 1478 341
rect 1462 322 1465 338
rect 1518 332 1521 358
rect 1526 352 1529 358
rect 1486 272 1489 318
rect 1494 312 1497 318
rect 1514 278 1518 281
rect 1526 272 1529 338
rect 1534 282 1537 448
rect 1542 342 1545 458
rect 1542 292 1545 328
rect 1498 268 1502 271
rect 1470 262 1473 268
rect 1534 262 1537 278
rect 1550 272 1553 498
rect 1558 492 1561 518
rect 1574 492 1577 548
rect 1598 542 1601 548
rect 1590 482 1593 538
rect 1606 532 1609 538
rect 1598 492 1601 518
rect 1566 472 1569 478
rect 1582 462 1585 468
rect 1590 462 1593 478
rect 1606 472 1609 478
rect 1614 462 1617 548
rect 1642 538 1646 541
rect 1622 492 1625 528
rect 1654 492 1657 638
rect 1662 562 1665 568
rect 1670 542 1673 648
rect 1686 642 1689 658
rect 1718 652 1721 668
rect 1742 662 1745 918
rect 1750 852 1753 1058
rect 1758 1022 1761 1078
rect 1774 1062 1777 1088
rect 1810 1078 1814 1081
rect 1822 1072 1825 1078
rect 1838 1072 1841 1168
rect 1890 1158 1894 1161
rect 1846 1142 1849 1158
rect 1854 1152 1857 1158
rect 1878 1152 1881 1158
rect 1874 1138 1878 1141
rect 1866 1128 1870 1131
rect 1846 1102 1849 1118
rect 1858 1078 1862 1081
rect 1786 1068 1790 1071
rect 1810 1068 1814 1071
rect 1870 1062 1873 1088
rect 1878 1072 1881 1098
rect 1894 1092 1897 1128
rect 1902 1122 1905 1148
rect 1942 1132 1945 1178
rect 1958 1142 1961 1268
rect 1966 1232 1969 1348
rect 1974 1332 1977 1418
rect 1982 1382 1985 1388
rect 1990 1342 1993 1348
rect 1998 1332 2001 1428
rect 2038 1402 2041 1458
rect 2058 1448 2062 1451
rect 2034 1388 2038 1391
rect 2006 1352 2009 1358
rect 2022 1352 2025 1358
rect 2046 1352 2049 1378
rect 2054 1362 2057 1448
rect 2070 1392 2073 1468
rect 2062 1352 2065 1358
rect 2054 1342 2057 1348
rect 2078 1332 2081 1528
rect 2094 1452 2097 1538
rect 2090 1448 2094 1451
rect 1990 1282 1993 1328
rect 2078 1312 2081 1328
rect 2014 1272 2017 1278
rect 2030 1272 2033 1308
rect 2070 1292 2073 1298
rect 2094 1292 2097 1418
rect 2102 1392 2105 1538
rect 2134 1532 2137 1548
rect 2158 1542 2161 1548
rect 2174 1532 2177 1638
rect 2310 1631 2313 1650
rect 2194 1568 2198 1571
rect 2182 1552 2185 1558
rect 2214 1552 2217 1608
rect 2222 1561 2225 1618
rect 2266 1568 2270 1571
rect 2222 1558 2230 1561
rect 2186 1528 2190 1531
rect 2134 1492 2137 1518
rect 2230 1492 2233 1558
rect 2286 1552 2289 1598
rect 2298 1558 2302 1561
rect 2250 1548 2254 1551
rect 2258 1538 2262 1541
rect 2262 1522 2265 1528
rect 2214 1472 2217 1478
rect 2230 1472 2233 1478
rect 2118 1462 2121 1468
rect 2302 1462 2305 1468
rect 2110 1452 2113 1458
rect 2130 1428 2134 1431
rect 2114 1378 2118 1381
rect 2102 1352 2105 1358
rect 2102 1322 2105 1348
rect 2158 1322 2161 1348
rect 2214 1342 2217 1438
rect 2262 1431 2265 1450
rect 2262 1362 2265 1388
rect 2270 1352 2273 1458
rect 2310 1452 2313 1458
rect 2318 1451 2321 1518
rect 2334 1502 2337 1538
rect 2350 1522 2353 1668
rect 2366 1662 2369 1668
rect 2358 1562 2361 1618
rect 2346 1518 2350 1521
rect 2334 1472 2337 1498
rect 2374 1492 2377 1538
rect 2326 1462 2329 1468
rect 2334 1462 2337 1468
rect 2358 1452 2361 1458
rect 2318 1448 2326 1451
rect 2286 1352 2289 1378
rect 2310 1362 2313 1428
rect 2298 1358 2302 1361
rect 2298 1348 2302 1351
rect 2286 1342 2289 1348
rect 2318 1342 2321 1378
rect 2342 1362 2345 1388
rect 2358 1382 2361 1388
rect 2326 1352 2329 1358
rect 2338 1348 2342 1351
rect 2374 1342 2377 1458
rect 2382 1422 2385 1688
rect 2486 1682 2489 1768
rect 2526 1752 2529 1818
rect 2534 1752 2537 1758
rect 2502 1692 2505 1728
rect 2394 1678 2398 1681
rect 2402 1658 2405 1661
rect 2502 1652 2505 1668
rect 2542 1662 2545 1858
rect 2654 1822 2657 1848
rect 2662 1822 2665 1858
rect 2686 1852 2689 1928
rect 2694 1872 2697 2138
rect 2710 2122 2713 2128
rect 2702 2092 2705 2118
rect 2734 2092 2737 2148
rect 2750 2112 2753 2268
rect 2802 2258 2806 2261
rect 2782 2231 2785 2250
rect 2822 2222 2825 2268
rect 2886 2262 2889 2268
rect 2842 2218 2846 2221
rect 2854 2152 2857 2258
rect 2870 2162 2873 2188
rect 2822 2142 2825 2148
rect 2894 2142 2897 2178
rect 2910 2162 2913 2188
rect 2926 2152 2929 2248
rect 2982 2202 2985 2338
rect 3030 2332 3033 2408
rect 3046 2352 3049 2378
rect 3054 2362 3057 2528
rect 3062 2512 3065 2518
rect 3070 2462 3073 2548
rect 3102 2522 3105 2538
rect 3126 2502 3129 2548
rect 3158 2542 3161 2548
rect 3138 2538 3142 2541
rect 3166 2532 3169 2538
rect 3086 2482 3089 2488
rect 3078 2472 3081 2478
rect 3094 2472 3097 2488
rect 3158 2482 3161 2528
rect 3110 2472 3113 2478
rect 3158 2472 3161 2478
rect 3166 2472 3169 2478
rect 3130 2468 3134 2471
rect 3070 2452 3073 2458
rect 3118 2442 3121 2458
rect 3142 2452 3145 2458
rect 3166 2452 3169 2458
rect 3134 2442 3137 2448
rect 3094 2352 3097 2368
rect 3118 2352 3121 2438
rect 3166 2432 3169 2448
rect 3174 2442 3177 2638
rect 3182 2632 3185 2668
rect 3218 2658 3222 2661
rect 3210 2648 3214 2651
rect 3182 2622 3185 2628
rect 3182 2542 3185 2618
rect 3198 2562 3201 2648
rect 3230 2642 3233 2668
rect 3238 2642 3241 2658
rect 3238 2592 3241 2638
rect 3246 2632 3249 2668
rect 3262 2642 3265 2668
rect 3278 2662 3281 2668
rect 3310 2662 3313 2668
rect 3366 2662 3369 2678
rect 3414 2662 3417 2668
rect 3518 2662 3521 2748
rect 3526 2712 3529 2738
rect 3542 2731 3545 2758
rect 3566 2752 3569 2758
rect 3550 2742 3553 2748
rect 3570 2738 3574 2741
rect 3586 2738 3590 2741
rect 3542 2728 3553 2731
rect 3534 2672 3537 2718
rect 3330 2658 3334 2661
rect 3250 2558 3254 2561
rect 3274 2558 3281 2561
rect 3190 2542 3193 2548
rect 3182 2492 3185 2538
rect 3198 2492 3201 2558
rect 3278 2552 3281 2558
rect 3234 2548 3238 2551
rect 3266 2548 3270 2551
rect 3206 2532 3209 2538
rect 3214 2522 3217 2548
rect 3294 2541 3297 2648
rect 3310 2562 3313 2578
rect 3326 2572 3329 2618
rect 3342 2582 3345 2658
rect 3330 2548 3334 2551
rect 3342 2542 3345 2548
rect 3290 2538 3297 2541
rect 3306 2538 3310 2541
rect 3214 2512 3217 2518
rect 3186 2478 3190 2481
rect 3214 2472 3217 2508
rect 3230 2492 3233 2538
rect 3250 2528 3254 2531
rect 3278 2502 3281 2538
rect 3294 2532 3297 2538
rect 3318 2522 3321 2538
rect 3246 2492 3249 2498
rect 3286 2492 3289 2518
rect 3318 2502 3321 2518
rect 3314 2488 3318 2491
rect 3222 2472 3225 2488
rect 3206 2462 3209 2468
rect 3254 2462 3257 2468
rect 3270 2462 3273 2478
rect 3214 2451 3217 2458
rect 3210 2448 3217 2451
rect 3246 2452 3249 2458
rect 3278 2452 3281 2478
rect 3294 2462 3297 2468
rect 3302 2462 3305 2478
rect 3318 2462 3321 2468
rect 3334 2452 3337 2528
rect 3350 2481 3353 2538
rect 3358 2492 3361 2518
rect 3350 2478 3361 2481
rect 3358 2462 3361 2478
rect 3366 2472 3369 2518
rect 3374 2472 3377 2628
rect 3382 2622 3385 2650
rect 3534 2642 3537 2668
rect 3542 2652 3545 2658
rect 3518 2622 3521 2638
rect 3472 2603 3474 2607
rect 3478 2603 3481 2607
rect 3485 2603 3488 2607
rect 3446 2532 3449 2598
rect 3510 2562 3513 2588
rect 3462 2542 3465 2548
rect 3414 2472 3417 2498
rect 3426 2478 3454 2481
rect 3378 2468 3382 2471
rect 3434 2468 3438 2471
rect 3366 2462 3369 2468
rect 3446 2462 3449 2468
rect 3486 2462 3489 2488
rect 3498 2478 3502 2481
rect 3494 2462 3497 2468
rect 3346 2458 3350 2461
rect 3418 2458 3422 2461
rect 3338 2448 3342 2451
rect 3146 2428 3150 2431
rect 3142 2392 3145 2418
rect 3166 2382 3169 2428
rect 3182 2372 3185 2378
rect 3190 2362 3193 2448
rect 3258 2438 3262 2441
rect 3398 2422 3401 2458
rect 3466 2448 3470 2451
rect 3406 2392 3409 2418
rect 3472 2403 3474 2407
rect 3478 2403 3481 2407
rect 3485 2403 3488 2407
rect 3162 2358 3166 2361
rect 3058 2348 3062 2351
rect 3178 2348 3182 2351
rect 3226 2348 3230 2351
rect 3070 2332 3073 2348
rect 3086 2342 3089 2348
rect 3130 2338 3134 2341
rect 3002 2328 3006 2331
rect 3078 2322 3081 2338
rect 3158 2332 3161 2348
rect 3190 2312 3193 2338
rect 3078 2262 3081 2268
rect 2994 2258 2998 2261
rect 2990 2222 2993 2248
rect 3034 2238 3038 2241
rect 3118 2232 3121 2278
rect 3134 2272 3137 2278
rect 3182 2262 3185 2278
rect 3198 2272 3201 2348
rect 3238 2342 3241 2368
rect 3502 2360 3505 2379
rect 3294 2352 3297 2358
rect 3266 2348 3270 2351
rect 3254 2342 3257 2348
rect 3206 2332 3209 2338
rect 3226 2328 3230 2331
rect 3214 2322 3217 2328
rect 3206 2302 3209 2318
rect 3206 2262 3209 2298
rect 3222 2271 3225 2328
rect 3218 2268 3225 2271
rect 3230 2272 3233 2318
rect 3262 2312 3265 2348
rect 3302 2342 3305 2348
rect 3310 2342 3313 2348
rect 3326 2342 3329 2358
rect 3282 2338 3286 2341
rect 3270 2332 3273 2338
rect 3334 2332 3337 2358
rect 3354 2348 3358 2351
rect 3282 2328 3286 2331
rect 3270 2312 3273 2328
rect 3302 2272 3305 2308
rect 3326 2272 3329 2328
rect 3334 2272 3337 2318
rect 3342 2312 3345 2338
rect 3358 2332 3361 2338
rect 3370 2318 3374 2321
rect 3342 2292 3345 2308
rect 3406 2302 3409 2348
rect 3310 2268 3318 2271
rect 3226 2258 3230 2261
rect 2958 2152 2961 2188
rect 2906 2138 2910 2141
rect 2806 2122 2809 2128
rect 2910 2122 2913 2128
rect 2734 2072 2737 2088
rect 2742 2072 2745 2108
rect 2838 2092 2841 2108
rect 2774 2072 2777 2078
rect 2798 2072 2801 2078
rect 2830 2072 2833 2078
rect 2714 2068 2718 2071
rect 2838 2062 2841 2078
rect 2862 2072 2865 2098
rect 2870 2082 2873 2088
rect 2894 2072 2897 2108
rect 2902 2072 2905 2098
rect 2910 2062 2913 2088
rect 2926 2082 2929 2148
rect 2982 2142 2985 2198
rect 2994 2168 2998 2171
rect 2938 2138 2942 2141
rect 2952 2103 2954 2107
rect 2958 2103 2961 2107
rect 2965 2103 2968 2107
rect 2850 2058 2854 2061
rect 2890 2058 2894 2061
rect 2922 2058 2926 2061
rect 2710 2052 2713 2058
rect 2726 2052 2729 2058
rect 2742 2022 2745 2058
rect 2762 2048 2766 2051
rect 2778 2048 2782 2051
rect 2750 2042 2753 2048
rect 2790 2042 2793 2048
rect 2798 2032 2801 2058
rect 2806 2042 2809 2048
rect 2822 2012 2825 2048
rect 2910 2042 2913 2058
rect 2926 2012 2929 2048
rect 2934 2002 2937 2068
rect 2846 1992 2849 1998
rect 2814 1962 2817 1988
rect 2942 1972 2945 2018
rect 2950 1992 2953 2068
rect 2818 1948 2822 1951
rect 2766 1942 2769 1948
rect 2886 1942 2889 1948
rect 2942 1942 2945 1948
rect 2974 1942 2977 2018
rect 2750 1922 2753 1928
rect 2714 1888 2718 1891
rect 2694 1862 2697 1868
rect 2726 1862 2729 1908
rect 2734 1862 2737 1868
rect 2706 1858 2710 1861
rect 2714 1848 2718 1851
rect 2586 1758 2590 1761
rect 2606 1752 2609 1788
rect 2654 1752 2657 1758
rect 2554 1738 2558 1741
rect 2610 1738 2614 1741
rect 2566 1722 2569 1738
rect 2574 1682 2577 1708
rect 2582 1692 2585 1738
rect 2630 1722 2633 1748
rect 2590 1672 2593 1678
rect 2622 1672 2625 1718
rect 2630 1662 2633 1718
rect 2602 1658 2606 1661
rect 2614 1652 2617 1658
rect 2630 1652 2633 1658
rect 2638 1652 2641 1658
rect 2602 1648 2606 1651
rect 2550 1622 2553 1648
rect 2440 1603 2442 1607
rect 2446 1603 2449 1607
rect 2453 1603 2456 1607
rect 2534 1592 2537 1598
rect 2470 1560 2473 1579
rect 2622 1571 2625 1628
rect 2646 1622 2649 1748
rect 2662 1742 2665 1818
rect 2686 1762 2689 1848
rect 2742 1842 2745 1878
rect 2790 1862 2793 1898
rect 2870 1892 2873 1928
rect 2798 1862 2801 1868
rect 2814 1862 2817 1868
rect 2882 1858 2886 1861
rect 2670 1722 2673 1728
rect 2686 1692 2689 1718
rect 2654 1672 2657 1678
rect 2686 1672 2689 1688
rect 2694 1682 2697 1838
rect 2758 1822 2761 1858
rect 2774 1842 2777 1848
rect 2702 1722 2705 1748
rect 2710 1742 2713 1758
rect 2734 1752 2737 1758
rect 2750 1742 2753 1818
rect 2758 1762 2761 1818
rect 2790 1762 2793 1858
rect 2806 1852 2809 1858
rect 2798 1762 2801 1838
rect 2814 1772 2817 1858
rect 2846 1792 2849 1818
rect 2878 1792 2881 1798
rect 2862 1762 2865 1768
rect 2826 1758 2830 1761
rect 2854 1758 2862 1761
rect 2826 1748 2830 1751
rect 2742 1732 2745 1738
rect 2766 1732 2769 1738
rect 2774 1732 2777 1738
rect 2782 1732 2785 1748
rect 2794 1738 2798 1741
rect 2714 1728 2718 1731
rect 2758 1702 2761 1718
rect 2806 1702 2809 1738
rect 2702 1692 2705 1698
rect 2662 1642 2665 1648
rect 2678 1622 2681 1658
rect 2678 1612 2681 1618
rect 2694 1602 2697 1678
rect 2750 1672 2753 1688
rect 2710 1652 2713 1658
rect 2718 1652 2721 1658
rect 2606 1568 2625 1571
rect 2606 1562 2609 1568
rect 2590 1558 2598 1561
rect 2550 1552 2553 1558
rect 2590 1552 2593 1558
rect 2614 1552 2617 1558
rect 2622 1552 2625 1568
rect 2718 1562 2721 1598
rect 2726 1562 2729 1658
rect 2734 1582 2737 1658
rect 2742 1632 2745 1668
rect 2766 1662 2769 1688
rect 2782 1682 2785 1688
rect 2806 1662 2809 1678
rect 2814 1672 2817 1748
rect 2754 1658 2758 1661
rect 2822 1652 2825 1748
rect 2838 1732 2841 1738
rect 2854 1732 2857 1758
rect 2878 1752 2881 1778
rect 2838 1702 2841 1728
rect 2862 1692 2865 1698
rect 2830 1682 2833 1688
rect 2870 1672 2873 1708
rect 2886 1692 2889 1738
rect 2918 1712 2921 1718
rect 2846 1662 2849 1668
rect 2830 1642 2833 1648
rect 2846 1642 2849 1658
rect 2886 1562 2889 1618
rect 2638 1552 2641 1558
rect 2562 1548 2566 1551
rect 2674 1548 2678 1551
rect 2438 1542 2441 1548
rect 2422 1532 2425 1538
rect 2486 1532 2489 1548
rect 2574 1542 2577 1548
rect 2510 1522 2513 1538
rect 2410 1488 2414 1491
rect 2422 1472 2425 1518
rect 2510 1482 2513 1518
rect 2394 1468 2398 1471
rect 2458 1468 2462 1471
rect 2482 1468 2485 1471
rect 2422 1462 2425 1468
rect 2526 1462 2529 1528
rect 2558 1502 2561 1538
rect 2590 1532 2593 1538
rect 2598 1522 2601 1548
rect 2654 1542 2657 1548
rect 2630 1522 2633 1538
rect 2670 1532 2673 1548
rect 2686 1542 2689 1558
rect 2642 1528 2646 1531
rect 2654 1502 2657 1528
rect 2686 1502 2689 1528
rect 2566 1482 2569 1488
rect 2654 1472 2657 1498
rect 2694 1491 2697 1518
rect 2686 1488 2697 1491
rect 2710 1492 2713 1548
rect 2718 1512 2721 1558
rect 2734 1552 2737 1558
rect 2826 1548 2830 1551
rect 2750 1542 2753 1548
rect 2782 1542 2785 1548
rect 2886 1542 2889 1548
rect 2742 1522 2745 1538
rect 2786 1528 2790 1531
rect 2686 1472 2689 1488
rect 2694 1472 2697 1478
rect 2674 1468 2678 1471
rect 2582 1462 2585 1468
rect 2634 1458 2638 1461
rect 2702 1461 2705 1478
rect 2734 1472 2737 1478
rect 2698 1458 2705 1461
rect 2398 1452 2401 1458
rect 2478 1452 2481 1458
rect 2418 1448 2422 1451
rect 2398 1362 2401 1448
rect 2438 1432 2441 1448
rect 2434 1418 2438 1421
rect 2440 1403 2442 1407
rect 2446 1403 2449 1407
rect 2453 1403 2456 1407
rect 2438 1362 2441 1388
rect 2386 1348 2390 1351
rect 2402 1348 2406 1351
rect 2198 1322 2201 1328
rect 2062 1282 2065 1288
rect 2190 1272 2193 1278
rect 2206 1272 2209 1278
rect 2026 1268 2030 1271
rect 2074 1268 2078 1271
rect 2286 1271 2289 1278
rect 2286 1268 2294 1271
rect 1990 1262 1993 1268
rect 2010 1258 2014 1261
rect 1982 1252 1985 1258
rect 1966 1158 1974 1161
rect 1986 1158 1990 1161
rect 1966 1152 1969 1158
rect 1998 1152 2001 1258
rect 2054 1222 2057 1268
rect 2062 1252 2065 1258
rect 2094 1192 2097 1248
rect 2106 1238 2110 1241
rect 2150 1202 2153 1258
rect 2238 1222 2241 1250
rect 2278 1242 2281 1268
rect 2290 1258 2294 1261
rect 2302 1222 2305 1238
rect 2322 1228 2326 1231
rect 2150 1160 2153 1179
rect 2166 1152 2169 1198
rect 1978 1148 1982 1151
rect 2118 1142 2121 1148
rect 1998 1132 2001 1138
rect 2014 1132 2017 1138
rect 1946 1128 1950 1131
rect 1918 1092 1921 1128
rect 2102 1122 2105 1128
rect 2018 1118 2022 1121
rect 1928 1103 1930 1107
rect 1934 1103 1937 1107
rect 1941 1103 1944 1107
rect 1950 1102 1953 1118
rect 2022 1092 2025 1108
rect 2062 1082 2065 1088
rect 1906 1078 1910 1081
rect 1978 1078 1982 1081
rect 2026 1078 2030 1081
rect 1930 1068 1934 1071
rect 1966 1071 1969 1078
rect 2094 1072 2097 1098
rect 1966 1068 1990 1071
rect 2106 1068 2110 1071
rect 1810 1058 1817 1061
rect 1782 1051 1785 1058
rect 1774 1048 1785 1051
rect 1774 1042 1777 1048
rect 1782 982 1785 1028
rect 1806 992 1809 1038
rect 1814 1012 1817 1058
rect 1774 962 1777 978
rect 1822 962 1825 1048
rect 1758 952 1761 958
rect 1758 892 1761 938
rect 1774 922 1777 958
rect 1794 948 1798 951
rect 1830 951 1833 1058
rect 1850 1048 1854 1051
rect 1878 1051 1881 1058
rect 1870 1048 1881 1051
rect 1870 1042 1873 1048
rect 1850 958 1854 961
rect 1862 952 1865 1008
rect 1902 992 1905 1058
rect 1910 1012 1913 1068
rect 1954 1058 1958 1061
rect 1942 992 1945 1058
rect 1990 1042 1993 1058
rect 2006 1022 2009 1058
rect 2026 1048 2030 1051
rect 1954 1018 1958 1021
rect 2038 982 2041 1018
rect 2046 1012 2049 1058
rect 2078 1052 2081 1068
rect 2118 1062 2121 1098
rect 2130 1078 2134 1081
rect 1994 978 1998 981
rect 1882 958 1886 961
rect 1982 952 1985 958
rect 2054 952 2057 958
rect 2078 952 2081 1048
rect 1822 948 1833 951
rect 1850 948 1854 951
rect 1874 948 1878 951
rect 1898 948 1902 951
rect 1930 948 1934 951
rect 1962 948 1966 951
rect 2034 948 2038 951
rect 1794 938 1798 941
rect 1806 932 1809 948
rect 1758 862 1761 878
rect 1766 862 1769 868
rect 1774 852 1777 918
rect 1782 872 1785 878
rect 1806 872 1809 878
rect 1822 872 1825 948
rect 1830 932 1833 938
rect 1878 932 1881 938
rect 1790 862 1793 868
rect 1798 842 1801 868
rect 1806 842 1809 858
rect 1806 792 1809 828
rect 1766 762 1769 768
rect 1786 758 1790 761
rect 1802 748 1806 751
rect 1814 751 1817 868
rect 1830 862 1833 878
rect 1838 872 1841 918
rect 1846 862 1849 868
rect 1898 858 1901 861
rect 1870 852 1873 858
rect 1822 792 1825 838
rect 1910 832 1913 938
rect 1922 928 1926 931
rect 1958 922 1961 928
rect 1974 922 1977 948
rect 2018 938 2022 941
rect 1928 903 1930 907
rect 1934 903 1937 907
rect 1941 903 1944 907
rect 1982 882 1985 888
rect 1998 872 2001 888
rect 2070 882 2073 948
rect 2094 941 2097 1058
rect 2126 992 2129 1018
rect 2102 952 2105 978
rect 2134 972 2137 1068
rect 2150 1062 2153 1118
rect 2166 1082 2169 1148
rect 2174 1082 2177 1198
rect 2194 1188 2198 1191
rect 2234 1158 2238 1161
rect 2254 1152 2257 1218
rect 2302 1202 2305 1218
rect 2350 1212 2353 1338
rect 2374 1332 2377 1338
rect 2430 1332 2433 1348
rect 2402 1328 2406 1331
rect 2406 1272 2409 1278
rect 2422 1272 2425 1278
rect 2462 1262 2465 1398
rect 2510 1392 2513 1418
rect 2526 1402 2529 1458
rect 2630 1422 2633 1448
rect 2470 1352 2473 1388
rect 2482 1378 2489 1381
rect 2498 1378 2502 1381
rect 2478 1342 2481 1378
rect 2486 1352 2489 1378
rect 2498 1348 2502 1351
rect 2510 1342 2513 1388
rect 2526 1342 2529 1358
rect 2550 1352 2553 1388
rect 2558 1341 2561 1378
rect 2566 1352 2569 1398
rect 2586 1358 2590 1361
rect 2574 1352 2577 1358
rect 2558 1338 2566 1341
rect 2470 1222 2473 1248
rect 2440 1203 2442 1207
rect 2446 1203 2449 1207
rect 2453 1203 2456 1207
rect 2270 1162 2273 1168
rect 2262 1152 2265 1158
rect 2194 1148 2198 1151
rect 2218 1148 2222 1151
rect 2282 1148 2286 1151
rect 2306 1148 2310 1151
rect 2190 1122 2193 1148
rect 2318 1142 2321 1158
rect 2206 1122 2209 1128
rect 2142 1052 2145 1058
rect 2142 992 2145 1008
rect 2114 948 2118 951
rect 2150 942 2153 1018
rect 2182 972 2185 1018
rect 2214 1012 2217 1138
rect 2238 1122 2241 1128
rect 2246 1122 2249 1138
rect 2286 1132 2289 1138
rect 2306 1128 2310 1131
rect 2338 1128 2342 1131
rect 2390 1122 2393 1148
rect 2430 1132 2433 1168
rect 2478 1152 2481 1258
rect 2486 1232 2489 1338
rect 2518 1282 2521 1288
rect 2510 1262 2513 1268
rect 2494 1162 2497 1188
rect 2526 1152 2529 1328
rect 2537 1258 2542 1261
rect 2574 1232 2577 1348
rect 2598 1332 2601 1348
rect 2614 1282 2617 1388
rect 2622 1352 2625 1358
rect 2630 1352 2633 1378
rect 2622 1322 2625 1328
rect 2638 1312 2641 1458
rect 2654 1452 2657 1458
rect 2710 1422 2713 1448
rect 2718 1412 2721 1468
rect 2726 1462 2729 1468
rect 2742 1462 2745 1518
rect 2870 1512 2873 1528
rect 2926 1512 2929 1928
rect 2952 1903 2954 1907
rect 2958 1903 2961 1907
rect 2965 1903 2968 1907
rect 2982 1902 2985 2138
rect 3078 2132 3081 2198
rect 3126 2160 3129 2179
rect 3134 2152 3137 2258
rect 3166 2231 3169 2250
rect 3238 2232 3241 2258
rect 3246 2242 3249 2268
rect 3258 2258 3262 2261
rect 3258 2248 3262 2251
rect 3230 2182 3233 2188
rect 3094 2132 3097 2138
rect 3078 2101 3081 2128
rect 3078 2098 3089 2101
rect 3086 2082 3089 2098
rect 2994 2058 2998 2061
rect 2990 1962 2993 1988
rect 3006 1982 3009 2018
rect 3014 1952 3017 2078
rect 3102 2072 3105 2078
rect 3134 2062 3137 2148
rect 3166 2142 3169 2148
rect 3182 2142 3185 2168
rect 3238 2152 3241 2168
rect 3194 2148 3198 2151
rect 3250 2148 3254 2151
rect 3206 2132 3209 2148
rect 3238 2142 3241 2148
rect 3262 2142 3265 2178
rect 3270 2152 3273 2188
rect 3278 2182 3281 2218
rect 3286 2162 3289 2258
rect 3294 2252 3297 2258
rect 3302 2222 3305 2268
rect 3310 2211 3313 2268
rect 3318 2242 3321 2248
rect 3326 2242 3329 2258
rect 3302 2208 3313 2211
rect 3334 2212 3337 2268
rect 3358 2262 3361 2298
rect 3390 2262 3393 2268
rect 3398 2262 3401 2298
rect 3414 2282 3417 2348
rect 3470 2342 3473 2358
rect 3510 2352 3513 2548
rect 3526 2472 3529 2478
rect 3542 2472 3545 2648
rect 3550 2632 3553 2728
rect 3590 2722 3593 2728
rect 3582 2702 3585 2718
rect 3598 2712 3601 2858
rect 3618 2848 3622 2851
rect 3630 2832 3633 2878
rect 3658 2858 3662 2861
rect 3646 2851 3649 2858
rect 3678 2852 3681 2858
rect 3646 2848 3657 2851
rect 3646 2752 3649 2808
rect 3654 2772 3657 2848
rect 3666 2838 3670 2841
rect 3686 2762 3689 2918
rect 3702 2892 3705 2928
rect 3710 2892 3713 2908
rect 3718 2902 3721 2918
rect 3710 2872 3713 2888
rect 3742 2878 3745 2948
rect 3762 2928 3766 2931
rect 3782 2892 3785 2958
rect 3846 2952 3849 3078
rect 3862 3042 3865 3068
rect 3886 3062 3889 3078
rect 3970 3068 3974 3071
rect 4082 3068 4086 3071
rect 3874 3058 3878 3061
rect 3902 3052 3905 3058
rect 3890 3038 3894 3041
rect 3878 3002 3881 3018
rect 3790 2892 3793 2948
rect 3854 2942 3857 2978
rect 3886 2952 3889 3018
rect 3902 3002 3905 3048
rect 3910 3022 3913 3068
rect 3926 3062 3929 3068
rect 3950 3052 3953 3058
rect 3930 3048 3934 3051
rect 3958 3022 3961 3068
rect 3958 2962 3961 2998
rect 3898 2958 3902 2961
rect 3946 2958 3950 2961
rect 3958 2942 3961 2958
rect 3926 2932 3929 2938
rect 3842 2928 3846 2931
rect 3766 2882 3769 2888
rect 3698 2868 3702 2871
rect 3770 2858 3774 2861
rect 3782 2852 3785 2868
rect 3806 2862 3809 2868
rect 3798 2852 3801 2858
rect 3814 2852 3817 2928
rect 3854 2892 3857 2928
rect 3886 2882 3889 2888
rect 3862 2872 3865 2878
rect 3910 2872 3913 2878
rect 3842 2858 3846 2861
rect 3854 2852 3857 2868
rect 3886 2862 3889 2868
rect 3838 2832 3841 2838
rect 3878 2832 3881 2848
rect 3886 2842 3889 2858
rect 3894 2842 3897 2858
rect 3910 2842 3913 2848
rect 3702 2762 3705 2818
rect 3742 2812 3745 2818
rect 3662 2752 3665 2758
rect 3746 2748 3750 2751
rect 3646 2742 3649 2748
rect 3582 2682 3585 2688
rect 3558 2662 3561 2668
rect 3566 2662 3569 2678
rect 3578 2668 3582 2671
rect 3598 2662 3601 2708
rect 3606 2672 3609 2708
rect 3614 2682 3617 2688
rect 3578 2648 3582 2651
rect 3606 2622 3609 2668
rect 3614 2662 3617 2668
rect 3630 2622 3633 2718
rect 3646 2692 3649 2728
rect 3654 2722 3657 2738
rect 3734 2732 3737 2748
rect 3758 2732 3761 2738
rect 3774 2732 3777 2808
rect 3794 2768 3798 2771
rect 3782 2752 3785 2758
rect 3798 2752 3801 2758
rect 3806 2741 3809 2748
rect 3802 2738 3809 2741
rect 3714 2728 3718 2731
rect 3698 2718 3702 2721
rect 3678 2672 3681 2698
rect 3702 2672 3705 2688
rect 3710 2672 3713 2698
rect 3718 2661 3721 2718
rect 3750 2662 3753 2718
rect 3774 2682 3777 2728
rect 3802 2688 3806 2691
rect 3790 2672 3793 2678
rect 3814 2672 3817 2808
rect 3838 2762 3841 2828
rect 3830 2758 3838 2761
rect 3830 2742 3833 2758
rect 3854 2752 3857 2828
rect 3918 2812 3921 2918
rect 3926 2872 3929 2918
rect 3966 2892 3969 3068
rect 4038 3062 4041 3068
rect 4102 3062 4105 3068
rect 3994 3058 3998 3061
rect 4010 3058 4014 3061
rect 4058 3058 4062 3061
rect 4114 3058 4118 3061
rect 3982 2952 3985 2958
rect 3990 2922 3993 3048
rect 3998 3042 4001 3048
rect 4022 3042 4025 3058
rect 4038 3052 4041 3058
rect 4030 3042 4033 3048
rect 4102 3032 4105 3058
rect 4110 3042 4113 3048
rect 4126 3032 4129 3038
rect 4046 3002 4049 3018
rect 3998 2982 4001 2988
rect 4054 2982 4057 3008
rect 4102 2992 4105 3028
rect 4038 2962 4041 2968
rect 4026 2948 4030 2951
rect 3976 2903 3978 2907
rect 3982 2903 3985 2907
rect 3989 2903 3992 2907
rect 3998 2902 4001 2948
rect 4006 2891 4009 2938
rect 4014 2932 4017 2948
rect 4054 2942 4057 2978
rect 4110 2972 4113 2978
rect 4118 2972 4121 3018
rect 4142 3012 4145 3068
rect 4150 3062 4153 3078
rect 4182 3062 4185 3078
rect 4202 3068 4206 3071
rect 4234 3068 4238 3071
rect 4250 3068 4254 3071
rect 4282 3068 4286 3071
rect 4306 3058 4310 3061
rect 4162 3048 4166 3051
rect 4174 3042 4177 3048
rect 4150 2972 4153 3018
rect 4166 2992 4169 3018
rect 4182 2972 4185 3058
rect 4190 3032 4193 3038
rect 4198 2982 4201 3018
rect 4138 2968 4142 2971
rect 4170 2968 4174 2971
rect 4042 2928 4046 2931
rect 4030 2912 4033 2928
rect 4062 2912 4065 2948
rect 4086 2942 4089 2968
rect 4154 2958 4158 2961
rect 4094 2952 4097 2958
rect 4102 2942 4105 2958
rect 4114 2948 4118 2951
rect 4154 2948 4158 2951
rect 4070 2932 4073 2938
rect 4150 2932 4153 2938
rect 4082 2928 4086 2931
rect 4134 2892 4137 2908
rect 4174 2902 4177 2958
rect 4190 2952 4193 2958
rect 4182 2912 4185 2948
rect 4198 2932 4201 2938
rect 4206 2932 4209 3048
rect 4214 2962 4217 2988
rect 4222 2922 4225 2958
rect 4230 2932 4233 3058
rect 4238 3022 4241 3058
rect 4270 3052 4273 3058
rect 4298 3048 4302 3051
rect 4314 3038 4318 3041
rect 4238 2942 4241 2998
rect 4246 2992 4249 3028
rect 4294 3022 4297 3028
rect 4262 3002 4265 3018
rect 4294 2992 4297 3008
rect 4326 2972 4329 3018
rect 4342 3002 4345 3018
rect 4370 2988 4374 2991
rect 4374 2972 4377 2978
rect 4266 2968 4273 2971
rect 4262 2962 4265 2968
rect 4258 2948 4262 2951
rect 4254 2922 4257 2928
rect 4166 2892 4169 2898
rect 4206 2892 4209 2918
rect 4230 2912 4233 2918
rect 4238 2892 4241 2918
rect 3998 2888 4009 2891
rect 3926 2862 3929 2868
rect 3934 2862 3937 2888
rect 3986 2878 3990 2881
rect 3942 2862 3945 2868
rect 3958 2862 3961 2868
rect 3966 2862 3969 2868
rect 3934 2832 3937 2858
rect 3946 2848 3950 2851
rect 3978 2848 3982 2851
rect 3842 2748 3846 2751
rect 3866 2748 3870 2751
rect 3834 2738 3838 2741
rect 3834 2728 3838 2731
rect 3854 2722 3857 2748
rect 3878 2741 3881 2768
rect 3874 2738 3881 2741
rect 3886 2742 3889 2778
rect 3946 2758 3950 2761
rect 3898 2748 3902 2751
rect 3986 2748 3990 2751
rect 3870 2681 3873 2728
rect 3902 2712 3905 2748
rect 3934 2732 3937 2748
rect 3866 2678 3873 2681
rect 3762 2668 3766 2671
rect 3806 2668 3814 2671
rect 3714 2658 3721 2661
rect 3738 2658 3742 2661
rect 3638 2612 3641 2658
rect 3662 2582 3665 2658
rect 3670 2652 3673 2658
rect 3774 2652 3777 2658
rect 3730 2648 3734 2651
rect 3766 2622 3769 2648
rect 3694 2602 3697 2618
rect 3550 2492 3553 2528
rect 3534 2462 3537 2468
rect 3558 2462 3561 2578
rect 3690 2558 3694 2561
rect 3586 2548 3590 2551
rect 3630 2542 3633 2558
rect 3614 2532 3617 2538
rect 3602 2528 3606 2531
rect 3570 2518 3574 2521
rect 3618 2518 3622 2521
rect 3566 2462 3569 2508
rect 3590 2462 3593 2488
rect 3610 2478 3614 2481
rect 3622 2462 3625 2468
rect 3630 2462 3633 2468
rect 3638 2462 3641 2538
rect 3646 2472 3649 2558
rect 3718 2551 3721 2558
rect 3782 2552 3785 2668
rect 3806 2652 3809 2668
rect 3822 2662 3825 2678
rect 3834 2668 3838 2671
rect 3870 2662 3873 2678
rect 3886 2672 3889 2678
rect 3894 2662 3897 2668
rect 3838 2632 3841 2648
rect 3790 2562 3793 2618
rect 3846 2612 3849 2618
rect 3854 2602 3857 2638
rect 3902 2632 3905 2708
rect 3918 2682 3921 2718
rect 3814 2552 3817 2558
rect 3714 2548 3721 2551
rect 3770 2548 3774 2551
rect 3654 2482 3657 2528
rect 3662 2502 3665 2538
rect 3670 2532 3673 2548
rect 3806 2542 3809 2548
rect 3682 2538 3686 2541
rect 3714 2538 3718 2541
rect 3762 2538 3766 2541
rect 3810 2538 3817 2541
rect 3694 2492 3697 2518
rect 3662 2482 3665 2488
rect 3694 2481 3697 2488
rect 3694 2478 3702 2481
rect 3710 2472 3713 2478
rect 3718 2472 3721 2488
rect 3690 2468 3694 2471
rect 3726 2462 3729 2508
rect 3742 2502 3745 2538
rect 3774 2532 3777 2538
rect 3754 2528 3758 2531
rect 3774 2472 3777 2508
rect 3782 2482 3785 2488
rect 3814 2462 3817 2538
rect 3842 2538 3846 2541
rect 3830 2532 3833 2538
rect 3522 2458 3526 2461
rect 3666 2458 3670 2461
rect 3770 2458 3774 2461
rect 3546 2448 3550 2451
rect 3550 2362 3553 2368
rect 3454 2292 3457 2328
rect 3502 2282 3505 2318
rect 3426 2278 3430 2281
rect 3422 2272 3425 2278
rect 3458 2268 3462 2271
rect 3406 2262 3409 2268
rect 3378 2258 3382 2261
rect 3450 2258 3454 2261
rect 3350 2252 3353 2258
rect 3382 2252 3385 2258
rect 3478 2252 3481 2258
rect 3486 2252 3489 2268
rect 3450 2228 3454 2231
rect 3302 2192 3305 2208
rect 3472 2203 3474 2207
rect 3478 2203 3481 2207
rect 3485 2203 3488 2207
rect 3422 2182 3425 2188
rect 3410 2178 3414 2181
rect 3374 2162 3377 2178
rect 3470 2152 3473 2168
rect 3494 2152 3497 2208
rect 3518 2192 3521 2348
rect 3558 2342 3561 2458
rect 3566 2272 3569 2448
rect 3606 2432 3609 2448
rect 3582 2372 3585 2418
rect 3630 2382 3633 2458
rect 3798 2432 3801 2448
rect 3658 2428 3662 2431
rect 3638 2362 3641 2388
rect 3822 2382 3825 2518
rect 3830 2481 3833 2528
rect 3838 2522 3841 2528
rect 3854 2492 3857 2598
rect 3886 2582 3889 2588
rect 3894 2562 3897 2618
rect 3910 2552 3913 2648
rect 3918 2641 3921 2668
rect 3934 2662 3937 2668
rect 3930 2648 3934 2651
rect 3942 2641 3945 2738
rect 3958 2662 3961 2748
rect 3978 2728 3982 2731
rect 3954 2658 3958 2661
rect 3966 2652 3969 2728
rect 3978 2718 3982 2721
rect 3976 2703 3978 2707
rect 3982 2703 3985 2707
rect 3989 2703 3992 2707
rect 3998 2692 4001 2888
rect 4030 2882 4033 2888
rect 4006 2872 4009 2878
rect 4014 2862 4017 2868
rect 4030 2852 4033 2868
rect 4022 2848 4030 2851
rect 4006 2742 4009 2778
rect 3998 2682 4001 2688
rect 3986 2678 3990 2681
rect 4006 2652 4009 2668
rect 3918 2638 3929 2641
rect 3942 2638 3950 2641
rect 3926 2592 3929 2638
rect 3958 2632 3961 2648
rect 3914 2548 3918 2551
rect 3870 2532 3873 2538
rect 3934 2532 3937 2628
rect 3950 2592 3953 2628
rect 3966 2602 3969 2648
rect 3970 2558 3974 2561
rect 3950 2542 3953 2548
rect 3942 2532 3945 2538
rect 3966 2532 3969 2548
rect 4006 2542 4009 2588
rect 4014 2582 4017 2658
rect 4022 2632 4025 2848
rect 4038 2842 4041 2888
rect 4242 2878 4246 2881
rect 4094 2872 4097 2878
rect 4126 2872 4129 2878
rect 4066 2868 4070 2871
rect 4138 2868 4142 2871
rect 4210 2868 4214 2871
rect 4242 2868 4246 2871
rect 4050 2858 4054 2861
rect 4114 2858 4118 2861
rect 4086 2852 4089 2858
rect 4090 2848 4097 2851
rect 4046 2832 4049 2838
rect 4030 2692 4033 2788
rect 4038 2762 4041 2798
rect 4038 2732 4041 2758
rect 4062 2752 4065 2758
rect 4078 2742 4081 2818
rect 4066 2738 4070 2741
rect 4082 2718 4086 2721
rect 4054 2712 4057 2718
rect 4046 2672 4049 2678
rect 4094 2672 4097 2848
rect 4126 2792 4129 2868
rect 4198 2862 4201 2868
rect 4254 2861 4257 2918
rect 4270 2872 4273 2968
rect 4346 2958 4350 2961
rect 4322 2948 4326 2951
rect 4278 2882 4281 2948
rect 4310 2942 4313 2948
rect 4286 2922 4289 2938
rect 4250 2858 4257 2861
rect 4110 2762 4113 2768
rect 4102 2692 4105 2748
rect 4126 2732 4129 2758
rect 4130 2728 4134 2731
rect 4034 2668 4038 2671
rect 4098 2668 4102 2671
rect 4118 2662 4121 2728
rect 4130 2718 4134 2721
rect 4142 2682 4145 2858
rect 4214 2852 4217 2858
rect 4150 2742 4153 2788
rect 4182 2752 4185 2818
rect 4246 2812 4249 2858
rect 4206 2792 4209 2808
rect 4166 2742 4169 2748
rect 4182 2702 4185 2718
rect 4190 2682 4193 2778
rect 4198 2762 4201 2768
rect 4214 2762 4217 2778
rect 4222 2762 4225 2798
rect 4242 2748 4246 2751
rect 4106 2648 4110 2651
rect 4038 2572 4041 2588
rect 4014 2542 4017 2548
rect 3862 2492 3865 2528
rect 3894 2512 3897 2518
rect 3890 2488 3894 2491
rect 3830 2478 3838 2481
rect 3918 2472 3921 2478
rect 3866 2468 3870 2471
rect 3846 2442 3849 2468
rect 3934 2462 3937 2528
rect 3990 2521 3993 2528
rect 3998 2521 4001 2528
rect 3990 2518 4001 2521
rect 3950 2462 3953 2518
rect 3976 2503 3978 2507
rect 3982 2503 3985 2507
rect 3989 2503 3992 2507
rect 3966 2482 3969 2488
rect 3982 2472 3985 2488
rect 3982 2462 3985 2468
rect 3926 2442 3929 2458
rect 3998 2442 4001 2518
rect 4014 2492 4017 2538
rect 4022 2532 4025 2558
rect 4030 2542 4033 2548
rect 4046 2541 4049 2648
rect 4118 2632 4121 2658
rect 4126 2642 4129 2668
rect 4134 2652 4137 2658
rect 4142 2652 4145 2658
rect 4166 2642 4169 2648
rect 4154 2638 4158 2641
rect 4078 2612 4081 2618
rect 4142 2592 4145 2618
rect 4054 2562 4057 2568
rect 4066 2558 4070 2561
rect 4046 2538 4054 2541
rect 4062 2532 4065 2538
rect 4022 2472 4025 2478
rect 4070 2462 4073 2548
rect 4078 2542 4081 2568
rect 4130 2548 4134 2551
rect 4138 2538 4142 2541
rect 4126 2532 4129 2538
rect 4078 2472 4081 2478
rect 4086 2462 4089 2518
rect 4082 2458 4086 2461
rect 4070 2452 4073 2458
rect 4018 2448 4022 2451
rect 3578 2358 3582 2361
rect 3574 2342 3577 2348
rect 3582 2281 3585 2338
rect 3590 2322 3593 2348
rect 3598 2342 3601 2358
rect 3634 2348 3638 2351
rect 3798 2342 3801 2368
rect 3818 2358 3822 2361
rect 3830 2351 3833 2418
rect 3902 2372 3905 2418
rect 3842 2358 3846 2361
rect 3830 2348 3838 2351
rect 3894 2342 3897 2358
rect 3902 2352 3905 2358
rect 3926 2342 3929 2368
rect 3998 2352 4001 2428
rect 4046 2352 4049 2418
rect 4054 2362 4057 2368
rect 4002 2348 4006 2351
rect 4050 2348 4057 2351
rect 4014 2342 4017 2348
rect 3818 2338 3822 2341
rect 3866 2338 3870 2341
rect 3618 2328 3622 2331
rect 3590 2292 3593 2298
rect 3606 2292 3609 2318
rect 3614 2282 3617 2318
rect 3686 2292 3689 2338
rect 3858 2328 3862 2331
rect 3582 2278 3593 2281
rect 3538 2268 3542 2271
rect 3566 2262 3569 2268
rect 3582 2262 3585 2268
rect 3590 2262 3593 2278
rect 3554 2258 3558 2261
rect 3526 2252 3529 2258
rect 3526 2232 3529 2238
rect 3542 2172 3545 2248
rect 3250 2138 3254 2141
rect 3166 2092 3169 2128
rect 3198 2092 3201 2118
rect 3214 2112 3217 2138
rect 3278 2132 3281 2148
rect 3286 2142 3289 2148
rect 3182 2072 3185 2078
rect 3206 2072 3209 2098
rect 3258 2088 3262 2091
rect 3230 2082 3233 2088
rect 3190 2062 3193 2068
rect 3198 2062 3201 2068
rect 3206 2062 3209 2068
rect 3214 2062 3217 2078
rect 3234 2068 3238 2071
rect 3246 2062 3249 2078
rect 3046 1952 3049 2058
rect 3170 2048 3174 2051
rect 3086 2022 3089 2048
rect 3054 1962 3057 2008
rect 2994 1948 2998 1951
rect 3062 1942 3065 1968
rect 3086 1962 3089 2018
rect 3070 1952 3073 1958
rect 3094 1942 3097 1978
rect 3134 1962 3137 2038
rect 3150 2022 3153 2048
rect 3106 1958 3110 1961
rect 3122 1948 3126 1951
rect 3130 1948 3134 1951
rect 3146 1948 3150 1951
rect 3026 1938 3030 1941
rect 3090 1938 3094 1941
rect 3058 1928 3062 1931
rect 3090 1928 3094 1931
rect 3102 1922 3105 1948
rect 3062 1892 3065 1918
rect 3118 1902 3121 1938
rect 3126 1922 3129 1938
rect 3158 1932 3161 1938
rect 3166 1932 3169 1958
rect 3182 1942 3185 1998
rect 3206 1971 3209 2058
rect 3246 2042 3249 2058
rect 3198 1968 3209 1971
rect 3198 1962 3201 1968
rect 3206 1952 3209 1958
rect 3214 1952 3217 1978
rect 3230 1952 3233 2028
rect 3254 1952 3257 2078
rect 3270 2072 3273 2088
rect 3278 2082 3281 2128
rect 3310 2102 3313 2148
rect 3342 2142 3345 2148
rect 3350 2142 3353 2148
rect 3298 2088 3302 2091
rect 3262 2052 3265 2058
rect 3278 2052 3281 2058
rect 3286 2002 3289 2068
rect 3310 2052 3313 2058
rect 3310 2002 3313 2048
rect 3294 1992 3297 1998
rect 3282 1978 3286 1981
rect 3194 1948 3198 1951
rect 3222 1942 3225 1948
rect 3310 1942 3313 1948
rect 3178 1938 3182 1941
rect 3258 1938 3262 1941
rect 3250 1928 3254 1931
rect 3178 1918 3182 1921
rect 2950 1872 2953 1878
rect 2974 1862 2977 1868
rect 2942 1672 2945 1858
rect 2998 1732 3001 1878
rect 3110 1872 3113 1888
rect 3118 1872 3121 1898
rect 3130 1888 3134 1891
rect 3142 1882 3145 1898
rect 3174 1892 3177 1898
rect 3090 1868 3094 1871
rect 3078 1862 3081 1868
rect 3102 1862 3105 1868
rect 3034 1818 3038 1821
rect 3046 1802 3049 1858
rect 3078 1852 3081 1858
rect 3086 1852 3089 1858
rect 3118 1822 3121 1858
rect 3142 1822 3145 1868
rect 3158 1862 3161 1888
rect 3206 1872 3209 1928
rect 3214 1872 3217 1888
rect 3234 1868 3238 1871
rect 3182 1862 3185 1868
rect 3198 1862 3201 1868
rect 3206 1862 3209 1868
rect 3246 1862 3249 1868
rect 3270 1862 3273 1938
rect 3318 1932 3321 2138
rect 3326 2122 3329 2128
rect 3334 2102 3337 2138
rect 3358 2122 3361 2148
rect 3370 2138 3374 2141
rect 3382 2112 3385 2148
rect 3414 2142 3417 2148
rect 3422 2142 3425 2148
rect 3390 2122 3393 2138
rect 3462 2132 3465 2138
rect 3410 2128 3414 2131
rect 3358 2082 3361 2108
rect 3382 2092 3385 2108
rect 3406 2082 3409 2128
rect 3338 2068 3342 2071
rect 3326 2062 3329 2068
rect 3326 1992 3329 2048
rect 3342 2042 3345 2058
rect 3358 2002 3361 2078
rect 3422 2072 3425 2078
rect 3438 2072 3441 2108
rect 3374 2062 3377 2068
rect 3406 2062 3409 2068
rect 3446 2062 3449 2128
rect 3502 2112 3505 2148
rect 3462 2092 3465 2098
rect 3490 2088 3494 2091
rect 3454 2072 3457 2078
rect 3470 2071 3473 2078
rect 3462 2068 3473 2071
rect 3450 2058 3454 2061
rect 3366 2052 3369 2058
rect 3390 1952 3393 2018
rect 3398 1992 3401 2058
rect 3410 2048 3414 2051
rect 3406 1952 3409 1958
rect 3346 1948 3350 1951
rect 3414 1942 3417 1978
rect 3430 1972 3433 2058
rect 3422 1952 3425 1958
rect 3446 1952 3449 2058
rect 3434 1948 3438 1951
rect 3462 1942 3465 2068
rect 3510 2062 3513 2158
rect 3526 2152 3529 2168
rect 3538 2138 3542 2141
rect 3522 2078 3526 2081
rect 3542 2072 3545 2088
rect 3522 2068 3526 2071
rect 3550 2062 3553 2118
rect 3558 2052 3561 2248
rect 3566 2232 3569 2258
rect 3578 2248 3582 2251
rect 3606 2242 3609 2268
rect 3590 2182 3593 2188
rect 3566 2152 3569 2158
rect 3566 2092 3569 2118
rect 3574 2092 3577 2148
rect 3582 2092 3585 2128
rect 3490 2048 3494 2051
rect 3472 2003 3474 2007
rect 3478 2003 3481 2007
rect 3485 2003 3488 2007
rect 3510 1962 3513 1968
rect 3518 1952 3521 2038
rect 3526 2032 3529 2038
rect 3526 1952 3529 1988
rect 3558 1962 3561 2048
rect 3574 2042 3577 2068
rect 3590 2052 3593 2168
rect 3606 2092 3609 2198
rect 3614 2192 3617 2278
rect 3678 2272 3681 2288
rect 3702 2281 3705 2328
rect 3894 2322 3897 2338
rect 4010 2328 4014 2331
rect 3954 2318 3958 2321
rect 3698 2278 3705 2281
rect 3666 2268 3670 2271
rect 3622 2241 3625 2258
rect 3630 2252 3633 2268
rect 3642 2258 3646 2261
rect 3654 2258 3662 2261
rect 3654 2252 3657 2258
rect 3638 2248 3646 2251
rect 3670 2251 3673 2258
rect 3666 2248 3673 2251
rect 3638 2241 3641 2248
rect 3622 2238 3641 2241
rect 3634 2148 3638 2151
rect 3614 2122 3617 2128
rect 3638 2112 3641 2138
rect 3626 2068 3630 2071
rect 3642 2068 3646 2071
rect 3586 2048 3590 2051
rect 3598 2051 3601 2068
rect 3642 2058 3646 2061
rect 3598 2048 3606 2051
rect 3606 2042 3609 2048
rect 3546 1958 3550 1961
rect 3554 1948 3558 1951
rect 3402 1938 3406 1941
rect 3458 1938 3462 1941
rect 3282 1928 3286 1931
rect 3278 1892 3281 1918
rect 3350 1912 3353 1938
rect 3358 1922 3361 1938
rect 3398 1932 3401 1938
rect 3438 1922 3441 1938
rect 3294 1862 3297 1898
rect 3154 1858 3158 1861
rect 3174 1852 3177 1858
rect 3186 1848 3190 1851
rect 3118 1792 3121 1818
rect 3046 1760 3049 1779
rect 3174 1762 3177 1848
rect 3182 1762 3185 1848
rect 3014 1742 3017 1758
rect 3106 1758 3110 1761
rect 3090 1748 3094 1751
rect 3122 1748 3126 1751
rect 2998 1712 3001 1728
rect 3054 1712 3057 1748
rect 3142 1742 3145 1758
rect 3182 1752 3185 1758
rect 3194 1748 3198 1751
rect 3150 1742 3153 1748
rect 3166 1742 3169 1748
rect 3078 1738 3086 1741
rect 2952 1703 2954 1707
rect 2958 1703 2961 1707
rect 2965 1703 2968 1707
rect 2974 1692 2977 1698
rect 2966 1622 2969 1668
rect 3030 1662 3033 1708
rect 3078 1702 3081 1738
rect 3118 1732 3121 1738
rect 3138 1728 3142 1731
rect 3070 1672 3073 1678
rect 3086 1672 3089 1708
rect 3166 1692 3169 1718
rect 3174 1702 3177 1738
rect 3190 1712 3193 1738
rect 3214 1732 3217 1778
rect 3198 1692 3201 1708
rect 3158 1662 3161 1668
rect 3206 1662 3209 1668
rect 3118 1622 3121 1650
rect 3126 1632 3129 1658
rect 2986 1618 2990 1621
rect 2934 1562 2937 1588
rect 3006 1560 3009 1579
rect 2942 1552 2945 1558
rect 2986 1548 2990 1551
rect 2774 1482 2777 1488
rect 2754 1468 2758 1471
rect 2734 1458 2742 1461
rect 2774 1461 2777 1478
rect 2782 1472 2785 1478
rect 2798 1462 2801 1488
rect 2834 1478 2838 1481
rect 2806 1472 2809 1478
rect 2846 1462 2849 1468
rect 2774 1458 2785 1461
rect 2734 1452 2737 1458
rect 2766 1452 2769 1458
rect 2746 1448 2750 1451
rect 2662 1352 2665 1358
rect 2654 1342 2657 1348
rect 2670 1342 2673 1408
rect 2682 1358 2686 1361
rect 2726 1352 2729 1378
rect 2734 1362 2737 1418
rect 2782 1352 2785 1458
rect 2826 1458 2830 1461
rect 2790 1452 2793 1458
rect 2814 1422 2817 1428
rect 2838 1422 2841 1428
rect 2854 1422 2857 1478
rect 2874 1458 2878 1461
rect 2898 1458 2901 1461
rect 2814 1372 2817 1418
rect 2790 1362 2793 1368
rect 2810 1358 2814 1361
rect 2830 1352 2833 1368
rect 2846 1362 2849 1398
rect 2878 1352 2881 1418
rect 2682 1348 2686 1351
rect 2810 1348 2814 1351
rect 2718 1342 2721 1348
rect 2774 1342 2777 1348
rect 2746 1338 2750 1341
rect 2650 1328 2654 1331
rect 2754 1328 2758 1331
rect 2782 1331 2785 1348
rect 2862 1342 2865 1348
rect 2886 1342 2889 1408
rect 2802 1338 2806 1341
rect 2774 1328 2785 1331
rect 2630 1272 2633 1288
rect 2670 1262 2673 1308
rect 2694 1261 2697 1278
rect 2702 1272 2705 1328
rect 2710 1272 2713 1328
rect 2722 1288 2726 1291
rect 2742 1272 2745 1278
rect 2766 1272 2769 1318
rect 2774 1282 2777 1328
rect 2730 1268 2734 1271
rect 2694 1258 2702 1261
rect 2662 1231 2665 1250
rect 2558 1152 2561 1218
rect 2570 1158 2574 1161
rect 2582 1152 2585 1158
rect 2554 1148 2558 1151
rect 2446 1122 2449 1138
rect 2526 1132 2529 1148
rect 2554 1138 2561 1141
rect 2294 1102 2297 1118
rect 2222 1062 2225 1078
rect 2262 1072 2265 1078
rect 2278 1052 2281 1068
rect 2318 1062 2321 1118
rect 2326 1082 2329 1118
rect 2350 1112 2353 1118
rect 2390 1108 2398 1111
rect 2310 1031 2313 1050
rect 2342 1021 2345 1098
rect 2390 1092 2393 1108
rect 2382 1082 2385 1088
rect 2350 1052 2353 1068
rect 2394 1058 2398 1061
rect 2342 1018 2353 1021
rect 2198 942 2201 948
rect 2094 938 2105 941
rect 2090 918 2094 921
rect 2102 892 2105 938
rect 2118 932 2121 938
rect 2134 932 2137 938
rect 2154 928 2158 931
rect 2118 882 2121 928
rect 2090 878 2094 881
rect 2098 878 2110 881
rect 1942 852 1945 858
rect 1814 748 1822 751
rect 1850 748 1854 751
rect 1766 682 1769 738
rect 1774 682 1777 688
rect 1782 682 1785 748
rect 1810 738 1814 741
rect 1750 672 1753 678
rect 1790 662 1793 688
rect 1730 658 1734 661
rect 1754 658 1758 661
rect 1678 552 1681 578
rect 1694 572 1697 638
rect 1726 592 1729 648
rect 1742 642 1745 648
rect 1694 562 1697 568
rect 1710 552 1713 568
rect 1742 552 1745 558
rect 1750 551 1753 658
rect 1766 592 1769 638
rect 1782 572 1785 618
rect 1794 568 1798 571
rect 1806 562 1809 618
rect 1814 592 1817 708
rect 1822 692 1825 748
rect 1838 722 1841 728
rect 1846 692 1849 698
rect 1826 688 1833 691
rect 1822 662 1825 678
rect 1746 548 1753 551
rect 1770 548 1774 551
rect 1562 448 1566 451
rect 1570 378 1574 381
rect 1566 352 1569 368
rect 1558 342 1561 348
rect 1582 341 1585 428
rect 1590 352 1593 358
rect 1582 338 1590 341
rect 1558 292 1561 338
rect 1566 272 1569 318
rect 1578 268 1582 271
rect 1498 258 1502 261
rect 1554 258 1558 261
rect 1462 252 1465 258
rect 1474 248 1478 251
rect 1530 248 1534 251
rect 1462 192 1465 248
rect 1458 158 1462 161
rect 1470 152 1473 228
rect 1482 218 1486 221
rect 1494 172 1497 178
rect 1534 162 1537 248
rect 1514 158 1518 161
rect 1494 152 1497 158
rect 1406 132 1409 148
rect 1526 142 1529 148
rect 1534 142 1537 148
rect 1550 142 1553 228
rect 1558 152 1561 258
rect 1566 142 1569 218
rect 1458 138 1462 141
rect 1574 141 1577 268
rect 1598 262 1601 308
rect 1606 292 1609 408
rect 1606 278 1614 281
rect 1594 248 1598 251
rect 1582 202 1585 218
rect 1586 178 1590 181
rect 1590 152 1593 158
rect 1598 152 1601 158
rect 1606 142 1609 278
rect 1622 272 1625 278
rect 1614 242 1617 268
rect 1630 182 1633 478
rect 1638 472 1641 488
rect 1638 282 1641 468
rect 1654 452 1657 478
rect 1686 472 1689 548
rect 1726 542 1729 548
rect 1710 492 1713 538
rect 1790 532 1793 558
rect 1810 548 1814 551
rect 1754 528 1758 531
rect 1778 528 1782 531
rect 1762 488 1766 491
rect 1750 482 1753 488
rect 1790 482 1793 528
rect 1662 458 1670 461
rect 1646 432 1649 438
rect 1646 392 1649 418
rect 1646 212 1649 318
rect 1662 232 1665 458
rect 1670 392 1673 398
rect 1694 372 1697 458
rect 1710 452 1713 478
rect 1742 462 1745 468
rect 1750 462 1753 478
rect 1766 462 1769 468
rect 1786 458 1790 461
rect 1774 452 1777 458
rect 1794 448 1798 451
rect 1718 411 1721 448
rect 1734 442 1737 448
rect 1710 408 1721 411
rect 1710 382 1713 408
rect 1774 391 1777 418
rect 1766 388 1777 391
rect 1694 332 1697 368
rect 1766 342 1769 388
rect 1750 332 1753 338
rect 1670 262 1673 288
rect 1710 282 1713 328
rect 1726 272 1729 288
rect 1798 282 1801 348
rect 1806 322 1809 528
rect 1814 472 1817 538
rect 1830 532 1833 688
rect 1822 522 1825 528
rect 1822 472 1825 478
rect 1830 472 1833 488
rect 1838 472 1841 658
rect 1846 552 1849 568
rect 1854 542 1857 718
rect 1862 662 1865 778
rect 1886 752 1889 758
rect 1934 752 1937 838
rect 1950 762 1953 808
rect 1982 792 1985 868
rect 2054 862 2057 868
rect 2030 831 2033 850
rect 2070 842 2073 858
rect 2046 792 2049 838
rect 2078 792 2081 798
rect 2014 762 2017 768
rect 2034 758 2038 761
rect 2066 758 2070 761
rect 1970 748 1974 751
rect 1986 748 1993 751
rect 2018 748 2022 751
rect 2042 748 2046 751
rect 1926 742 1929 748
rect 1894 732 1897 738
rect 1914 728 1918 731
rect 1870 712 1873 728
rect 1878 691 1881 718
rect 1870 688 1881 691
rect 1902 692 1905 718
rect 1910 712 1913 728
rect 1870 662 1873 688
rect 1878 678 1886 681
rect 1878 592 1881 678
rect 1898 658 1902 661
rect 1874 548 1878 551
rect 1886 551 1889 618
rect 1910 592 1913 678
rect 1918 592 1921 718
rect 1974 712 1977 738
rect 1966 708 1974 711
rect 1928 703 1930 707
rect 1934 703 1937 707
rect 1941 703 1944 707
rect 1942 662 1945 668
rect 1882 548 1889 551
rect 1898 548 1902 551
rect 1870 532 1873 548
rect 1878 532 1881 538
rect 1850 528 1854 531
rect 1866 458 1870 461
rect 1814 362 1817 388
rect 1782 262 1785 278
rect 1806 272 1809 318
rect 1814 292 1817 298
rect 1822 272 1825 308
rect 1830 272 1833 448
rect 1838 402 1841 458
rect 1854 412 1857 448
rect 1838 352 1841 378
rect 1846 352 1849 358
rect 1846 312 1849 338
rect 1818 268 1822 271
rect 1830 262 1833 268
rect 1794 258 1798 261
rect 1774 222 1777 248
rect 1782 232 1785 258
rect 1630 152 1633 178
rect 1618 148 1622 151
rect 1742 142 1745 198
rect 1782 152 1785 228
rect 1842 218 1846 221
rect 1854 192 1857 358
rect 1862 342 1865 448
rect 1790 162 1793 188
rect 1574 138 1582 141
rect 1618 138 1622 141
rect 1642 138 1645 141
rect 1406 92 1409 108
rect 1338 88 1342 91
rect 1326 72 1329 78
rect 1306 68 1311 71
rect 1310 62 1313 68
rect 1366 62 1369 88
rect 1398 72 1401 78
rect 1378 68 1382 71
rect 1142 52 1145 58
rect 1086 32 1089 38
rect 1182 31 1185 50
rect 1342 32 1345 38
rect 1398 22 1401 38
rect 1430 22 1433 38
rect 790 -22 801 -19
rect 886 -19 890 -18
rect 894 -19 897 18
rect 886 -22 897 -19
rect 958 -19 962 -18
rect 966 -19 969 18
rect 958 -22 969 -19
rect 982 -19 986 -18
rect 990 -19 993 18
rect 982 -22 993 -19
rect 1006 -18 1009 8
rect 1006 -22 1010 -18
rect 1070 -19 1074 -18
rect 1078 -19 1081 18
rect 1070 -22 1081 -19
rect 1198 -18 1201 8
rect 1198 -22 1202 -18
rect 1350 -19 1353 18
rect 1374 -18 1377 8
rect 1416 3 1418 7
rect 1422 3 1425 7
rect 1429 3 1432 7
rect 1438 -18 1441 128
rect 1446 62 1449 138
rect 1566 132 1569 138
rect 1726 132 1729 138
rect 1478 102 1481 118
rect 1598 92 1601 108
rect 1622 102 1625 118
rect 1726 102 1729 128
rect 1622 92 1625 98
rect 1518 82 1521 88
rect 1702 82 1705 98
rect 1502 72 1505 78
rect 1718 72 1721 78
rect 1662 62 1665 68
rect 1782 62 1785 148
rect 1830 142 1833 148
rect 1862 142 1865 278
rect 1870 262 1873 348
rect 1878 282 1881 468
rect 1894 462 1897 528
rect 1910 492 1913 578
rect 1934 572 1937 618
rect 1918 562 1921 568
rect 1934 552 1937 568
rect 1942 552 1945 588
rect 1958 552 1961 618
rect 1928 503 1930 507
rect 1934 503 1937 507
rect 1941 503 1944 507
rect 1950 502 1953 548
rect 1966 542 1969 708
rect 1978 678 1982 681
rect 1974 602 1977 658
rect 1974 552 1977 598
rect 1982 562 1985 618
rect 1990 601 1993 748
rect 1998 732 2001 738
rect 2006 722 2009 738
rect 1998 692 2001 718
rect 1990 598 1998 601
rect 1990 562 1993 568
rect 1998 552 2001 598
rect 1986 538 1990 541
rect 2014 532 2017 728
rect 2022 612 2025 748
rect 2086 742 2089 878
rect 2166 872 2169 938
rect 2238 932 2241 978
rect 2302 962 2305 988
rect 2326 952 2329 1008
rect 2342 942 2345 1008
rect 2350 942 2353 1018
rect 2358 1012 2361 1058
rect 2366 1052 2369 1058
rect 2358 952 2361 958
rect 2366 952 2369 998
rect 2338 938 2342 941
rect 2254 932 2257 938
rect 2346 928 2350 931
rect 2238 912 2241 928
rect 2166 862 2169 868
rect 2094 772 2097 858
rect 2206 782 2209 878
rect 2222 872 2225 878
rect 2294 862 2297 868
rect 2310 862 2313 898
rect 2366 872 2369 938
rect 2374 932 2377 1048
rect 2422 1042 2425 1078
rect 2438 1062 2441 1108
rect 2534 1102 2537 1138
rect 2542 1102 2545 1118
rect 2558 1092 2561 1138
rect 2582 1132 2585 1148
rect 2606 1132 2609 1218
rect 2614 1152 2617 1178
rect 2622 1172 2625 1178
rect 2678 1152 2681 1258
rect 2710 1222 2713 1268
rect 2754 1258 2758 1261
rect 2742 1251 2745 1258
rect 2742 1248 2750 1251
rect 2766 1160 2769 1179
rect 2774 1162 2777 1278
rect 2790 1272 2793 1318
rect 2814 1292 2817 1338
rect 2838 1331 2841 1338
rect 2854 1332 2857 1338
rect 2838 1328 2846 1331
rect 2898 1328 2902 1331
rect 2826 1278 2830 1281
rect 2806 1272 2809 1278
rect 2838 1272 2841 1328
rect 2790 1262 2793 1268
rect 2798 1262 2801 1268
rect 2870 1262 2873 1308
rect 2910 1282 2913 1508
rect 2952 1503 2954 1507
rect 2958 1503 2961 1507
rect 2965 1503 2968 1507
rect 2982 1482 2985 1518
rect 3038 1512 3041 1538
rect 3054 1522 3057 1528
rect 3102 1482 3105 1488
rect 3106 1468 3110 1471
rect 2998 1402 3001 1468
rect 3086 1462 3089 1468
rect 3126 1462 3129 1628
rect 3134 1592 3137 1648
rect 3182 1642 3185 1658
rect 3194 1648 3198 1651
rect 3134 1552 3137 1588
rect 3142 1562 3145 1588
rect 3182 1582 3185 1638
rect 3222 1612 3225 1858
rect 3238 1812 3241 1848
rect 3246 1762 3249 1858
rect 3246 1752 3249 1758
rect 3230 1742 3233 1748
rect 3238 1742 3241 1748
rect 3050 1458 3054 1461
rect 3090 1448 3094 1451
rect 3046 1422 3049 1448
rect 2966 1352 2969 1358
rect 2922 1348 2926 1351
rect 2950 1342 2953 1348
rect 2938 1338 2942 1341
rect 2634 1148 2637 1151
rect 2810 1148 2814 1151
rect 2614 1142 2617 1148
rect 2574 1092 2577 1128
rect 2462 1082 2465 1088
rect 2538 1078 2542 1081
rect 2546 1068 2550 1071
rect 2478 1062 2481 1068
rect 2558 1062 2561 1088
rect 2430 1042 2433 1058
rect 2382 932 2385 1038
rect 2438 1031 2441 1058
rect 2430 1028 2441 1031
rect 2390 932 2393 968
rect 2398 932 2401 1018
rect 2430 952 2433 1028
rect 2440 1003 2442 1007
rect 2446 1003 2449 1007
rect 2453 1003 2456 1007
rect 2478 962 2481 968
rect 2486 952 2489 1018
rect 2502 952 2505 958
rect 2518 952 2521 998
rect 2582 992 2585 1108
rect 2598 1082 2601 1118
rect 2606 1092 2609 1128
rect 2614 1092 2617 1128
rect 2638 1072 2641 1088
rect 2678 1082 2681 1148
rect 2718 1122 2721 1128
rect 2734 1122 2737 1138
rect 2822 1132 2825 1168
rect 2870 1162 2873 1198
rect 2910 1192 2913 1278
rect 2926 1272 2929 1338
rect 2966 1332 2969 1348
rect 2952 1303 2954 1307
rect 2958 1303 2961 1307
rect 2965 1303 2968 1307
rect 2990 1282 2993 1338
rect 2998 1252 3001 1358
rect 3018 1348 3022 1351
rect 3018 1338 3022 1341
rect 3022 1312 3025 1338
rect 3038 1322 3041 1328
rect 3010 1268 3014 1271
rect 2974 1222 2977 1248
rect 3018 1218 3022 1221
rect 2898 1168 2905 1171
rect 2902 1162 2905 1168
rect 2842 1158 2846 1161
rect 2854 1152 2857 1158
rect 2870 1152 2873 1158
rect 2878 1152 2881 1158
rect 2842 1148 2846 1151
rect 2894 1142 2897 1158
rect 2926 1152 2929 1188
rect 2934 1152 2937 1158
rect 2922 1148 2926 1151
rect 2654 1072 2657 1078
rect 2674 1068 2677 1071
rect 2718 1062 2721 1078
rect 2758 1072 2761 1078
rect 2774 1062 2777 1068
rect 2626 1058 2630 1061
rect 2598 992 2601 1058
rect 2474 948 2478 951
rect 2514 948 2518 951
rect 2406 942 2409 948
rect 2374 912 2377 918
rect 2382 892 2385 918
rect 2398 872 2401 918
rect 2422 872 2425 928
rect 2430 882 2433 948
rect 2446 932 2449 948
rect 2534 942 2537 948
rect 2542 942 2545 978
rect 2622 962 2625 968
rect 2630 962 2633 1058
rect 2654 1052 2657 1058
rect 2662 1052 2665 1058
rect 2550 952 2553 958
rect 2670 952 2673 998
rect 2686 992 2689 1048
rect 2806 1031 2809 1050
rect 2734 962 2737 1008
rect 2746 968 2750 971
rect 2758 962 2761 978
rect 2790 962 2793 968
rect 2734 952 2737 958
rect 2814 952 2817 1118
rect 2822 1072 2825 1128
rect 2830 1102 2833 1138
rect 2862 1122 2865 1138
rect 2926 1122 2929 1138
rect 2950 1122 2953 1148
rect 2982 1142 2985 1178
rect 2990 1152 2993 1198
rect 3022 1162 3025 1198
rect 3006 1152 3009 1158
rect 2846 1082 2849 1118
rect 2894 1092 2897 1108
rect 2926 1102 2929 1118
rect 2934 1082 2937 1118
rect 2952 1103 2954 1107
rect 2958 1103 2961 1107
rect 2965 1103 2968 1107
rect 2890 1078 2894 1081
rect 2962 1078 2966 1081
rect 2846 952 2849 1078
rect 2862 1062 2865 1078
rect 2918 1072 2921 1078
rect 2946 1068 2950 1071
rect 2870 1062 2873 1068
rect 2854 992 2857 1018
rect 2866 958 2870 961
rect 2886 952 2889 1058
rect 2894 992 2897 1048
rect 2918 962 2921 1068
rect 2974 1062 2977 1138
rect 3006 1122 3009 1128
rect 3014 1122 3017 1138
rect 2990 1072 2993 1098
rect 2938 1058 2942 1061
rect 3002 1058 3006 1061
rect 2962 1048 2966 1051
rect 2926 972 2929 1048
rect 3010 1028 3014 1031
rect 2626 948 2630 951
rect 2770 948 2774 951
rect 2802 948 2806 951
rect 2662 942 2665 948
rect 2686 942 2689 948
rect 2514 938 2526 941
rect 2618 938 2622 941
rect 2746 938 2750 941
rect 2770 938 2777 941
rect 2446 892 2449 928
rect 2454 912 2457 938
rect 2354 868 2358 871
rect 2410 868 2414 871
rect 2410 858 2414 861
rect 2302 852 2305 858
rect 2438 852 2441 858
rect 2254 822 2257 850
rect 2342 842 2345 848
rect 2362 838 2366 841
rect 2158 742 2161 778
rect 2222 762 2225 788
rect 2302 752 2305 778
rect 2250 748 2254 751
rect 2222 742 2225 748
rect 2294 742 2297 748
rect 2038 722 2041 738
rect 2078 682 2081 728
rect 2086 702 2089 738
rect 2158 732 2161 738
rect 2174 732 2177 738
rect 2134 682 2137 698
rect 2182 682 2185 698
rect 2078 621 2081 678
rect 2094 672 2097 678
rect 2070 618 2081 621
rect 2038 562 2041 568
rect 2022 542 2025 548
rect 2046 542 2049 548
rect 2054 532 2057 538
rect 2018 528 2022 531
rect 1950 472 1953 498
rect 2006 492 2009 518
rect 2030 512 2033 518
rect 1894 452 1897 458
rect 1950 362 1953 468
rect 1982 342 1985 358
rect 1990 342 1993 478
rect 2006 442 2009 468
rect 2038 462 2041 488
rect 2026 388 2030 391
rect 2006 352 2009 358
rect 1938 338 1942 341
rect 1886 332 1889 338
rect 1928 303 1930 307
rect 1934 303 1937 307
rect 1941 303 1944 307
rect 1926 282 1929 288
rect 1990 272 1993 318
rect 1886 232 1889 258
rect 1942 232 1945 268
rect 1998 262 2001 328
rect 2014 292 2017 338
rect 2038 332 2041 458
rect 2054 422 2057 448
rect 2070 422 2073 618
rect 2086 502 2089 548
rect 2094 492 2097 658
rect 2118 552 2121 558
rect 2134 532 2137 678
rect 2190 672 2193 688
rect 2214 678 2230 681
rect 2198 662 2201 668
rect 2214 662 2217 678
rect 2222 662 2225 668
rect 2162 658 2166 661
rect 2230 652 2233 668
rect 2142 622 2145 648
rect 2106 518 2110 521
rect 2134 472 2137 518
rect 2142 472 2145 588
rect 2150 552 2153 558
rect 2158 552 2161 608
rect 2166 592 2169 598
rect 2162 538 2166 541
rect 2090 468 2094 471
rect 2078 452 2081 468
rect 2114 448 2118 451
rect 2126 442 2129 448
rect 2090 418 2094 421
rect 2102 412 2105 418
rect 2070 332 2073 348
rect 2110 342 2113 418
rect 2134 392 2137 458
rect 2142 452 2145 468
rect 2158 452 2161 478
rect 2174 472 2177 648
rect 2230 642 2233 648
rect 2210 638 2214 641
rect 2246 582 2249 728
rect 2254 642 2257 668
rect 2262 642 2265 648
rect 2262 632 2265 638
rect 2182 562 2185 568
rect 2222 562 2225 568
rect 2206 552 2209 558
rect 2218 548 2222 551
rect 2210 538 2214 541
rect 2186 528 2190 531
rect 2146 438 2150 441
rect 2166 352 2169 438
rect 2174 362 2177 388
rect 2198 342 2201 498
rect 2206 352 2209 528
rect 2238 512 2241 558
rect 2246 542 2249 578
rect 2270 561 2273 738
rect 2278 722 2281 728
rect 2286 722 2289 728
rect 2286 672 2289 688
rect 2278 612 2281 658
rect 2286 652 2289 658
rect 2294 652 2297 678
rect 2278 562 2281 568
rect 2270 558 2278 561
rect 2254 542 2257 548
rect 2294 542 2297 548
rect 2262 522 2265 538
rect 2302 532 2305 678
rect 2310 672 2313 818
rect 2326 762 2329 818
rect 2366 792 2369 828
rect 2390 762 2393 848
rect 2454 822 2457 908
rect 2470 872 2473 938
rect 2494 932 2497 938
rect 2510 922 2513 928
rect 2478 882 2481 888
rect 2486 872 2489 888
rect 2494 862 2497 878
rect 2502 872 2505 908
rect 2526 882 2529 938
rect 2590 922 2593 938
rect 2598 932 2601 938
rect 2534 882 2537 918
rect 2566 902 2569 918
rect 2590 902 2593 918
rect 2606 892 2609 918
rect 2614 912 2617 938
rect 2646 922 2649 928
rect 2598 882 2601 888
rect 2586 878 2590 881
rect 2518 872 2521 878
rect 2578 868 2582 871
rect 2550 862 2553 868
rect 2514 858 2518 861
rect 2462 852 2465 858
rect 2558 852 2561 858
rect 2566 842 2569 848
rect 2318 702 2321 718
rect 2326 692 2329 758
rect 2354 748 2358 751
rect 2402 748 2406 751
rect 2414 742 2417 818
rect 2440 803 2442 807
rect 2446 803 2449 807
rect 2453 803 2456 807
rect 2462 802 2465 828
rect 2354 738 2358 741
rect 2402 738 2406 741
rect 2318 681 2321 688
rect 2318 678 2329 681
rect 2326 662 2329 678
rect 2334 662 2337 718
rect 2366 692 2369 708
rect 2354 678 2358 681
rect 2314 658 2318 661
rect 2350 652 2353 658
rect 2374 652 2377 688
rect 2338 648 2342 651
rect 2350 642 2353 648
rect 2254 482 2257 488
rect 2270 472 2273 478
rect 2302 431 2305 450
rect 2242 388 2246 391
rect 2286 362 2289 398
rect 2310 362 2313 638
rect 2318 542 2321 588
rect 2350 572 2353 618
rect 2326 552 2329 558
rect 2350 542 2353 568
rect 2318 462 2321 538
rect 2338 528 2342 531
rect 2358 522 2361 548
rect 2374 541 2377 648
rect 2382 602 2385 738
rect 2390 682 2393 738
rect 2398 672 2401 718
rect 2422 712 2425 748
rect 2390 572 2393 658
rect 2406 562 2409 578
rect 2394 558 2398 561
rect 2386 548 2390 551
rect 2374 538 2382 541
rect 2338 518 2342 521
rect 2362 518 2369 521
rect 2366 472 2369 518
rect 2374 472 2377 518
rect 2422 502 2425 598
rect 2422 492 2425 498
rect 2390 472 2393 478
rect 2406 462 2409 468
rect 2354 458 2358 461
rect 2366 451 2369 458
rect 2362 448 2369 451
rect 2394 448 2398 451
rect 2282 358 2286 361
rect 2254 352 2257 358
rect 2274 348 2278 351
rect 2282 348 2286 351
rect 2110 332 2113 338
rect 2126 312 2129 338
rect 2206 302 2209 348
rect 2242 338 2246 341
rect 1974 222 1977 250
rect 2014 222 2017 288
rect 2026 268 2030 271
rect 2066 268 2070 271
rect 2038 262 2041 268
rect 1894 142 1897 208
rect 2018 178 2022 181
rect 1926 152 1929 158
rect 1906 148 1910 151
rect 1950 142 1953 158
rect 1958 152 1961 158
rect 1898 138 1902 141
rect 1798 92 1801 128
rect 1814 122 1817 138
rect 1918 102 1921 138
rect 1928 103 1930 107
rect 1934 103 1937 107
rect 1941 103 1944 107
rect 1794 88 1798 91
rect 1878 82 1881 88
rect 1894 62 1897 68
rect 1966 62 1969 138
rect 1974 132 1977 148
rect 2022 142 2025 148
rect 2030 142 2033 258
rect 2042 228 2046 231
rect 2038 152 2041 158
rect 2054 152 2057 208
rect 2078 162 2081 298
rect 2086 282 2089 288
rect 2094 282 2097 288
rect 2126 272 2129 278
rect 2158 272 2161 298
rect 2222 292 2225 318
rect 2166 272 2169 288
rect 2086 268 2102 271
rect 2202 268 2206 271
rect 2086 252 2089 268
rect 2094 248 2102 251
rect 2086 162 2089 218
rect 2078 152 2081 158
rect 2066 148 2070 151
rect 1998 132 2001 138
rect 2006 122 2009 128
rect 2014 82 2017 128
rect 1986 68 1990 71
rect 2014 62 2017 68
rect 2030 62 2033 138
rect 2046 132 2049 148
rect 2086 142 2089 148
rect 2058 138 2062 141
rect 2094 122 2097 248
rect 2118 232 2121 258
rect 2134 222 2137 248
rect 2110 168 2126 171
rect 2142 171 2145 268
rect 2150 252 2153 258
rect 2158 241 2161 258
rect 2230 252 2233 328
rect 2262 322 2265 338
rect 2278 322 2281 338
rect 2238 271 2241 318
rect 2238 268 2246 271
rect 2258 268 2262 271
rect 2278 262 2281 298
rect 2294 292 2297 348
rect 2310 342 2313 358
rect 2318 352 2321 358
rect 2310 332 2313 338
rect 2326 292 2329 448
rect 2342 402 2345 448
rect 2334 352 2337 368
rect 2346 358 2350 361
rect 2366 352 2369 428
rect 2366 342 2369 348
rect 2338 338 2342 341
rect 2378 338 2382 341
rect 2358 332 2361 338
rect 2378 328 2382 331
rect 2390 322 2393 328
rect 2398 302 2401 338
rect 2382 292 2385 298
rect 2366 282 2369 288
rect 2310 272 2313 278
rect 2370 268 2374 271
rect 2154 238 2161 241
rect 2214 248 2222 251
rect 2174 202 2177 218
rect 2142 168 2153 171
rect 2110 161 2113 168
rect 2102 158 2113 161
rect 2102 152 2105 158
rect 2126 152 2129 158
rect 2142 152 2145 158
rect 2110 142 2113 148
rect 2118 142 2121 148
rect 2046 92 2049 118
rect 2142 92 2145 148
rect 2150 142 2153 168
rect 2174 152 2177 158
rect 2182 152 2185 228
rect 2190 152 2193 158
rect 2158 102 2161 118
rect 2174 92 2177 138
rect 2190 92 2193 148
rect 2198 142 2201 178
rect 2118 82 2121 88
rect 2194 78 2198 81
rect 2062 72 2065 78
rect 2150 72 2153 78
rect 2162 68 2166 71
rect 2054 62 2057 68
rect 2206 62 2209 148
rect 2214 142 2217 248
rect 2238 192 2241 228
rect 2226 188 2230 191
rect 2254 172 2257 258
rect 2282 248 2286 251
rect 2302 202 2305 268
rect 2382 262 2385 288
rect 2398 262 2401 298
rect 2406 292 2409 458
rect 2430 352 2433 778
rect 2442 758 2446 761
rect 2462 752 2465 798
rect 2494 762 2497 838
rect 2574 801 2577 838
rect 2566 798 2577 801
rect 2566 792 2569 798
rect 2478 752 2481 758
rect 2442 748 2446 751
rect 2514 748 2518 751
rect 2470 712 2473 738
rect 2502 732 2505 738
rect 2518 732 2521 738
rect 2486 702 2489 728
rect 2526 702 2529 748
rect 2558 742 2561 778
rect 2574 762 2577 768
rect 2582 752 2585 758
rect 2590 751 2593 868
rect 2606 812 2609 868
rect 2614 862 2617 898
rect 2662 892 2665 938
rect 2678 932 2681 938
rect 2734 931 2737 938
rect 2734 928 2745 931
rect 2710 922 2713 928
rect 2674 878 2678 881
rect 2622 872 2625 878
rect 2694 872 2697 878
rect 2710 872 2713 918
rect 2742 892 2745 928
rect 2774 892 2777 938
rect 2814 941 2817 948
rect 2814 938 2822 941
rect 2806 922 2809 938
rect 2826 928 2830 931
rect 2782 872 2785 878
rect 2790 872 2793 918
rect 2806 912 2809 918
rect 2814 912 2817 918
rect 2822 882 2825 898
rect 2822 872 2825 878
rect 2830 872 2833 908
rect 2838 902 2841 948
rect 2846 932 2849 938
rect 2870 932 2873 938
rect 2878 892 2881 948
rect 2666 868 2670 871
rect 2754 868 2758 871
rect 2766 862 2769 868
rect 2626 858 2630 861
rect 2794 858 2798 861
rect 2602 768 2606 771
rect 2602 758 2609 761
rect 2590 748 2601 751
rect 2598 742 2601 748
rect 2606 742 2609 758
rect 2630 752 2633 828
rect 2638 812 2641 858
rect 2654 852 2657 858
rect 2638 762 2641 768
rect 2618 738 2622 741
rect 2534 732 2537 738
rect 2558 732 2561 738
rect 2550 722 2553 728
rect 2542 682 2545 718
rect 2582 692 2585 738
rect 2598 712 2601 738
rect 2590 692 2593 708
rect 2606 702 2609 728
rect 2440 603 2442 607
rect 2446 603 2449 607
rect 2453 603 2456 607
rect 2442 588 2446 591
rect 2478 552 2481 608
rect 2486 602 2489 678
rect 2502 672 2505 678
rect 2614 672 2617 708
rect 2646 692 2649 848
rect 2662 802 2665 848
rect 2734 822 2737 858
rect 2806 852 2809 868
rect 2742 822 2745 848
rect 2782 842 2785 848
rect 2774 822 2777 828
rect 2678 812 2681 818
rect 2678 792 2681 798
rect 2658 768 2662 771
rect 2654 742 2657 748
rect 2670 742 2673 748
rect 2626 688 2630 691
rect 2502 612 2505 658
rect 2534 622 2537 650
rect 2478 542 2481 548
rect 2534 542 2537 598
rect 2574 592 2577 668
rect 2610 658 2614 661
rect 2630 652 2633 678
rect 2654 672 2657 728
rect 2670 682 2673 738
rect 2662 672 2665 678
rect 2666 658 2670 661
rect 2686 652 2689 808
rect 2774 782 2777 818
rect 2814 802 2817 868
rect 2838 862 2841 878
rect 2870 872 2873 878
rect 2894 872 2897 958
rect 2902 922 2905 938
rect 2914 928 2918 931
rect 2926 872 2929 898
rect 2934 872 2937 938
rect 3030 932 3033 1298
rect 3038 1262 3041 1318
rect 3046 1272 3049 1398
rect 3070 1362 3073 1448
rect 3142 1441 3145 1558
rect 3174 1552 3177 1558
rect 3166 1542 3169 1548
rect 3150 1532 3153 1538
rect 3182 1532 3185 1548
rect 3214 1542 3217 1548
rect 3158 1522 3161 1528
rect 3206 1482 3209 1528
rect 3222 1502 3225 1518
rect 3238 1502 3241 1738
rect 3254 1662 3257 1818
rect 3278 1812 3281 1848
rect 3310 1842 3313 1868
rect 3326 1852 3329 1858
rect 3330 1838 3334 1841
rect 3266 1778 3270 1781
rect 3278 1752 3281 1778
rect 3298 1758 3302 1761
rect 3350 1752 3353 1908
rect 3358 1812 3361 1918
rect 3446 1902 3449 1918
rect 3510 1912 3513 1948
rect 3526 1942 3529 1948
rect 3534 1942 3537 1948
rect 3542 1932 3545 1938
rect 3574 1922 3577 1928
rect 3582 1912 3585 2008
rect 3598 1952 3601 2018
rect 3622 1992 3625 2058
rect 3630 1992 3633 2038
rect 3654 2012 3657 2058
rect 3662 1992 3665 2228
rect 3694 2192 3697 2278
rect 3738 2268 3742 2271
rect 3702 2222 3705 2268
rect 3710 2262 3713 2268
rect 3718 2242 3721 2268
rect 3766 2262 3769 2308
rect 3782 2272 3785 2318
rect 3746 2258 3750 2261
rect 3786 2258 3790 2261
rect 3726 2242 3729 2248
rect 3702 2162 3705 2218
rect 3678 2072 3681 2158
rect 3706 2138 3710 2141
rect 3678 2062 3681 2068
rect 3686 1992 3689 2068
rect 3710 2062 3713 2098
rect 3718 2092 3721 2238
rect 3734 2172 3737 2248
rect 3758 2212 3761 2258
rect 3814 2242 3817 2318
rect 3822 2262 3825 2268
rect 3822 2232 3825 2248
rect 3774 2162 3777 2228
rect 3730 2158 3734 2161
rect 3754 2158 3758 2161
rect 3802 2158 3806 2161
rect 3750 2142 3753 2148
rect 3782 2142 3785 2148
rect 3806 2142 3809 2148
rect 3830 2142 3833 2318
rect 3854 2272 3857 2318
rect 3862 2272 3865 2278
rect 3842 2258 3846 2261
rect 3886 2261 3889 2318
rect 3918 2302 3921 2318
rect 3914 2278 3918 2281
rect 3934 2262 3937 2318
rect 3976 2303 3978 2307
rect 3982 2303 3985 2307
rect 3989 2303 3992 2307
rect 3942 2272 3945 2298
rect 4014 2282 4017 2328
rect 3986 2278 3990 2281
rect 4002 2278 4006 2281
rect 4018 2268 4030 2271
rect 4054 2262 4057 2348
rect 4070 2322 4073 2338
rect 4086 2292 4089 2318
rect 4086 2262 4089 2278
rect 4094 2272 4097 2438
rect 4102 2431 4105 2518
rect 4150 2501 4153 2598
rect 4158 2562 4161 2628
rect 4162 2558 4166 2561
rect 4174 2552 4177 2678
rect 4150 2498 4161 2501
rect 4150 2472 4153 2488
rect 4142 2468 4150 2471
rect 4134 2462 4137 2468
rect 4114 2458 4118 2461
rect 4102 2428 4113 2431
rect 4102 2372 4105 2418
rect 4110 2361 4113 2428
rect 4106 2358 4113 2361
rect 4118 2352 4121 2368
rect 4134 2352 4137 2358
rect 4118 2342 4121 2348
rect 4142 2272 4145 2468
rect 4158 2462 4161 2498
rect 4182 2492 4185 2668
rect 4190 2551 4193 2678
rect 4198 2562 4201 2748
rect 4206 2722 4209 2748
rect 4222 2742 4225 2748
rect 4242 2738 4246 2741
rect 4270 2732 4273 2748
rect 4258 2728 4262 2731
rect 4206 2708 4209 2718
rect 4254 2672 4257 2718
rect 4230 2652 4233 2658
rect 4190 2548 4201 2551
rect 4190 2492 4193 2538
rect 4182 2452 4185 2488
rect 4198 2472 4201 2548
rect 4214 2542 4217 2568
rect 4158 2442 4161 2448
rect 4174 2422 4177 2448
rect 4150 2362 4153 2368
rect 4158 2332 4161 2418
rect 4198 2392 4201 2468
rect 4206 2452 4209 2518
rect 4214 2461 4217 2538
rect 4222 2532 4225 2628
rect 4246 2582 4249 2668
rect 4262 2662 4265 2688
rect 4278 2672 4281 2848
rect 4286 2822 4289 2878
rect 4294 2862 4297 2898
rect 4310 2882 4313 2938
rect 4318 2922 4321 2928
rect 4318 2872 4321 2898
rect 4334 2872 4337 2958
rect 4346 2948 4350 2951
rect 4358 2941 4361 2958
rect 4366 2952 4369 2958
rect 4354 2938 4361 2941
rect 4286 2792 4289 2818
rect 4294 2771 4297 2858
rect 4318 2852 4321 2858
rect 4306 2848 4310 2851
rect 4286 2768 4297 2771
rect 4314 2768 4318 2771
rect 4286 2672 4289 2768
rect 4294 2758 4302 2761
rect 4334 2752 4337 2868
rect 4350 2862 4353 2938
rect 4362 2848 4366 2851
rect 4310 2742 4313 2748
rect 4382 2742 4385 2858
rect 4330 2738 4334 2741
rect 4294 2722 4297 2738
rect 4318 2691 4321 2718
rect 4318 2688 4326 2691
rect 4334 2672 4337 2728
rect 4350 2712 4353 2718
rect 4382 2702 4385 2738
rect 4390 2702 4393 3058
rect 4390 2672 4393 2678
rect 4278 2662 4281 2668
rect 4286 2662 4289 2668
rect 4342 2662 4345 2668
rect 4306 2658 4310 2661
rect 4282 2648 4286 2651
rect 4246 2552 4249 2578
rect 4234 2548 4238 2551
rect 4270 2542 4273 2578
rect 4342 2552 4345 2648
rect 4350 2562 4353 2618
rect 4318 2542 4321 2548
rect 4358 2532 4361 2618
rect 4370 2558 4374 2561
rect 4378 2538 4390 2541
rect 4230 2482 4233 2518
rect 4302 2472 4305 2518
rect 4318 2492 4321 2528
rect 4358 2491 4361 2518
rect 4374 2492 4377 2518
rect 4358 2488 4369 2491
rect 4358 2472 4361 2478
rect 4226 2468 4230 2471
rect 4330 2468 4334 2471
rect 4214 2458 4222 2461
rect 4182 2362 4185 2368
rect 4222 2362 4225 2418
rect 4238 2402 4241 2468
rect 4290 2458 4294 2461
rect 4354 2458 4358 2461
rect 4270 2452 4273 2458
rect 4234 2358 4238 2361
rect 4198 2352 4201 2358
rect 4186 2348 4193 2351
rect 4150 2292 4153 2318
rect 4158 2272 4161 2328
rect 4190 2292 4193 2348
rect 4202 2338 4206 2341
rect 4214 2312 4217 2348
rect 4222 2332 4225 2338
rect 4166 2262 4169 2278
rect 4174 2272 4177 2278
rect 3886 2258 3894 2261
rect 3938 2258 3942 2261
rect 4002 2258 4006 2261
rect 4018 2258 4022 2261
rect 4042 2258 4046 2261
rect 4170 2258 4177 2261
rect 3950 2252 3953 2258
rect 3958 2248 3966 2251
rect 3838 2242 3841 2248
rect 3846 2192 3849 2218
rect 3854 2172 3857 2248
rect 3878 2242 3881 2248
rect 3934 2242 3937 2248
rect 3838 2142 3841 2148
rect 3730 2138 3734 2141
rect 3758 2132 3761 2138
rect 3774 2132 3777 2138
rect 3854 2132 3857 2168
rect 3862 2132 3865 2198
rect 3886 2162 3889 2238
rect 3902 2202 3905 2238
rect 3914 2218 3918 2221
rect 3910 2192 3913 2208
rect 3950 2162 3953 2218
rect 3958 2202 3961 2248
rect 3958 2192 3961 2198
rect 3998 2192 4001 2258
rect 4030 2242 4033 2258
rect 4146 2248 4150 2251
rect 4062 2242 4065 2248
rect 4126 2242 4129 2248
rect 4030 2192 4033 2238
rect 3898 2148 3902 2151
rect 3834 2128 3838 2131
rect 3822 2122 3825 2128
rect 3726 2092 3729 2118
rect 3734 2082 3737 2118
rect 3766 2072 3769 2078
rect 3794 2068 3798 2071
rect 3718 2062 3721 2068
rect 3706 2058 3710 2061
rect 3754 2058 3758 2061
rect 3606 1952 3609 1958
rect 3622 1952 3625 1968
rect 3702 1962 3705 2048
rect 3758 2042 3761 2048
rect 3710 1992 3713 2038
rect 3766 1991 3769 2068
rect 3774 2052 3777 2058
rect 3782 2032 3785 2068
rect 3806 2062 3809 2098
rect 3830 2082 3833 2088
rect 3854 2082 3857 2118
rect 3870 2092 3873 2138
rect 3886 2132 3889 2138
rect 3846 2062 3849 2068
rect 3878 2062 3881 2098
rect 3918 2082 3921 2138
rect 3926 2132 3929 2148
rect 3966 2142 3969 2168
rect 4046 2161 4049 2218
rect 4150 2182 4153 2188
rect 4134 2162 4137 2178
rect 4166 2162 4169 2168
rect 4038 2158 4049 2161
rect 4082 2158 4086 2161
rect 3934 2082 3937 2088
rect 3894 2062 3897 2068
rect 3918 2062 3921 2068
rect 3814 2052 3817 2058
rect 3854 2022 3857 2058
rect 3910 2042 3913 2048
rect 3766 1988 3777 1991
rect 3762 1978 3766 1981
rect 3730 1948 3734 1951
rect 3590 1942 3593 1948
rect 3622 1942 3625 1948
rect 3630 1932 3633 1948
rect 3646 1932 3649 1948
rect 3694 1942 3697 1948
rect 3718 1942 3721 1948
rect 3674 1938 3678 1941
rect 3414 1872 3417 1878
rect 3430 1872 3433 1878
rect 3518 1862 3521 1898
rect 3538 1888 3542 1891
rect 3542 1872 3545 1878
rect 3558 1872 3561 1878
rect 3530 1868 3534 1871
rect 3554 1868 3558 1871
rect 3514 1858 3518 1861
rect 3374 1822 3377 1858
rect 3462 1831 3465 1850
rect 3362 1768 3366 1771
rect 3374 1762 3377 1778
rect 3366 1752 3369 1758
rect 3330 1748 3334 1751
rect 3262 1702 3265 1748
rect 3270 1742 3273 1748
rect 3278 1742 3281 1748
rect 3286 1712 3289 1748
rect 3294 1742 3297 1748
rect 3338 1738 3342 1741
rect 3310 1722 3313 1738
rect 3350 1732 3353 1748
rect 3334 1702 3337 1718
rect 3374 1712 3377 1718
rect 3254 1632 3257 1658
rect 3246 1552 3249 1558
rect 3254 1522 3257 1528
rect 3222 1472 3225 1478
rect 3142 1438 3153 1441
rect 3074 1358 3081 1361
rect 3054 1272 3057 1348
rect 3070 1292 3073 1318
rect 3050 1258 3054 1261
rect 3038 1202 3041 1258
rect 3070 1252 3073 1278
rect 3038 1162 3041 1168
rect 3058 1158 3062 1161
rect 3078 1161 3081 1358
rect 3086 1272 3089 1408
rect 3150 1332 3153 1438
rect 3166 1352 3169 1458
rect 3254 1422 3257 1450
rect 3214 1362 3217 1388
rect 3234 1358 3238 1361
rect 3262 1352 3265 1578
rect 3270 1562 3273 1608
rect 3294 1592 3297 1678
rect 3310 1672 3313 1698
rect 3382 1662 3385 1808
rect 3472 1803 3474 1807
rect 3478 1803 3481 1807
rect 3485 1803 3488 1807
rect 3390 1722 3393 1748
rect 3398 1742 3401 1748
rect 3406 1742 3409 1768
rect 3430 1752 3433 1768
rect 3454 1752 3457 1758
rect 3462 1742 3465 1748
rect 3426 1738 3430 1741
rect 3390 1682 3393 1718
rect 3406 1712 3409 1728
rect 3414 1692 3417 1698
rect 3414 1672 3417 1688
rect 3410 1658 3414 1661
rect 3342 1631 3345 1650
rect 3326 1582 3329 1588
rect 3270 1552 3273 1558
rect 3286 1552 3289 1578
rect 3310 1562 3313 1568
rect 3342 1562 3345 1568
rect 3298 1558 3302 1561
rect 3330 1558 3337 1561
rect 3334 1552 3337 1558
rect 3366 1552 3369 1558
rect 3374 1552 3377 1628
rect 3382 1612 3385 1658
rect 3382 1592 3385 1598
rect 3398 1572 3401 1618
rect 3414 1592 3417 1658
rect 3390 1568 3398 1571
rect 3378 1548 3382 1551
rect 3278 1532 3281 1538
rect 3334 1532 3337 1538
rect 3302 1522 3305 1528
rect 3350 1522 3353 1538
rect 3366 1532 3369 1538
rect 3374 1532 3377 1538
rect 3390 1511 3393 1568
rect 3398 1552 3401 1558
rect 3406 1542 3409 1578
rect 3414 1552 3417 1558
rect 3430 1552 3433 1738
rect 3438 1722 3441 1728
rect 3442 1688 3446 1691
rect 3442 1668 3446 1671
rect 3494 1662 3497 1678
rect 3450 1658 3454 1661
rect 3466 1648 3470 1651
rect 3438 1632 3441 1648
rect 3442 1578 3446 1581
rect 3462 1562 3465 1648
rect 3472 1603 3474 1607
rect 3478 1603 3481 1607
rect 3485 1603 3488 1607
rect 3502 1592 3505 1748
rect 3510 1742 3513 1748
rect 3470 1562 3473 1568
rect 3494 1552 3497 1588
rect 3510 1552 3513 1678
rect 3526 1672 3529 1868
rect 3582 1862 3585 1908
rect 3590 1872 3593 1928
rect 3622 1882 3625 1918
rect 3594 1868 3598 1871
rect 3622 1862 3625 1878
rect 3630 1868 3638 1871
rect 3554 1858 3558 1861
rect 3610 1858 3614 1861
rect 3598 1852 3601 1858
rect 3630 1852 3633 1868
rect 3646 1862 3649 1898
rect 3654 1861 3657 1928
rect 3678 1922 3681 1928
rect 3702 1912 3705 1928
rect 3726 1892 3729 1918
rect 3742 1892 3745 1918
rect 3706 1888 3710 1891
rect 3662 1878 3689 1881
rect 3706 1878 3710 1881
rect 3662 1872 3665 1878
rect 3686 1872 3689 1878
rect 3742 1872 3745 1878
rect 3670 1868 3678 1871
rect 3654 1858 3665 1861
rect 3534 1752 3537 1818
rect 3550 1742 3553 1798
rect 3602 1768 3606 1771
rect 3618 1758 3622 1761
rect 3614 1752 3617 1758
rect 3586 1748 3590 1751
rect 3546 1718 3550 1721
rect 3542 1692 3545 1708
rect 3558 1672 3561 1738
rect 3614 1732 3617 1738
rect 3586 1728 3590 1731
rect 3566 1712 3569 1718
rect 3622 1712 3625 1748
rect 3630 1692 3633 1848
rect 3654 1791 3657 1848
rect 3662 1822 3665 1858
rect 3670 1842 3673 1868
rect 3690 1858 3694 1861
rect 3678 1852 3681 1858
rect 3718 1832 3721 1868
rect 3758 1862 3761 1868
rect 3766 1862 3769 1878
rect 3774 1872 3777 1988
rect 3782 1942 3785 2018
rect 3846 1932 3849 2008
rect 3910 1962 3913 1988
rect 3918 1972 3921 2018
rect 3862 1942 3865 1948
rect 3806 1882 3809 1888
rect 3878 1882 3881 1908
rect 3790 1872 3793 1878
rect 3822 1862 3825 1868
rect 3862 1862 3865 1878
rect 3894 1872 3897 1918
rect 3902 1912 3905 1948
rect 3934 1942 3937 2078
rect 3942 2062 3945 2118
rect 4014 2112 4017 2148
rect 4038 2141 4041 2158
rect 4050 2148 4054 2151
rect 4062 2142 4065 2158
rect 4098 2148 4102 2151
rect 4038 2138 4054 2141
rect 4106 2138 4110 2141
rect 4122 2138 4126 2141
rect 4134 2132 4137 2158
rect 4174 2152 4177 2258
rect 4182 2252 4185 2278
rect 4198 2272 4201 2278
rect 4214 2272 4217 2278
rect 4222 2272 4225 2318
rect 4246 2272 4249 2418
rect 4254 2352 4257 2398
rect 4286 2362 4289 2408
rect 4294 2392 4297 2448
rect 4318 2442 4321 2448
rect 4258 2348 4262 2351
rect 4314 2348 4321 2351
rect 4306 2338 4310 2341
rect 4254 2312 4257 2338
rect 4254 2282 4257 2288
rect 4190 2162 4193 2268
rect 4198 2172 4201 2258
rect 4190 2152 4193 2158
rect 4198 2152 4201 2168
rect 4154 2148 4158 2151
rect 4146 2138 4150 2141
rect 4174 2132 4177 2148
rect 4066 2128 4070 2131
rect 4082 2128 4094 2131
rect 3976 2103 3978 2107
rect 3982 2103 3985 2107
rect 3989 2103 3992 2107
rect 4002 2068 4006 2071
rect 4014 2052 4017 2108
rect 4070 2082 4073 2088
rect 4078 2082 4081 2098
rect 4026 2068 4030 2071
rect 4054 2062 4057 2068
rect 4046 2042 4049 2048
rect 3950 2012 3953 2018
rect 4010 1958 4014 1961
rect 4018 1958 4025 1961
rect 3958 1952 3961 1958
rect 3954 1948 3958 1951
rect 4014 1942 4017 1948
rect 3970 1938 3974 1941
rect 3934 1932 3937 1938
rect 4022 1932 4025 1958
rect 4074 1948 4078 1951
rect 4086 1942 4089 2118
rect 4118 2072 4121 2078
rect 4102 2062 4105 2068
rect 4126 2062 4129 2118
rect 4110 2052 4113 2058
rect 4094 2032 4097 2038
rect 4102 1961 4105 2018
rect 4118 1992 4121 2038
rect 4102 1958 4113 1961
rect 4094 1952 4097 1958
rect 4038 1932 4041 1938
rect 4070 1932 4073 1938
rect 3786 1858 3790 1861
rect 3914 1858 3918 1861
rect 3734 1852 3737 1858
rect 3774 1842 3777 1848
rect 3830 1842 3833 1858
rect 3934 1852 3937 1898
rect 3942 1872 3945 1918
rect 3958 1882 3961 1918
rect 3976 1903 3978 1907
rect 3982 1903 3985 1907
rect 3989 1903 3992 1907
rect 4006 1892 4009 1918
rect 3998 1872 4001 1878
rect 3970 1858 3974 1861
rect 3994 1858 3998 1861
rect 3898 1848 3902 1851
rect 3650 1788 3657 1791
rect 3638 1762 3641 1768
rect 3646 1762 3649 1788
rect 3726 1782 3729 1818
rect 3742 1792 3745 1818
rect 3662 1752 3665 1778
rect 3678 1742 3681 1758
rect 3602 1678 3606 1681
rect 3646 1672 3649 1708
rect 3654 1681 3657 1738
rect 3686 1692 3689 1748
rect 3702 1742 3705 1758
rect 3734 1752 3737 1758
rect 3726 1742 3729 1748
rect 3750 1742 3753 1808
rect 3758 1802 3761 1818
rect 3774 1792 3777 1838
rect 3758 1782 3761 1788
rect 3766 1742 3769 1748
rect 3778 1738 3782 1741
rect 3718 1702 3721 1718
rect 3686 1682 3689 1688
rect 3654 1678 3665 1681
rect 3530 1668 3534 1671
rect 3610 1668 3614 1671
rect 3634 1668 3641 1671
rect 3518 1661 3521 1668
rect 3518 1658 3526 1661
rect 3518 1642 3521 1648
rect 3422 1548 3430 1551
rect 3422 1542 3425 1548
rect 3430 1538 3438 1541
rect 3430 1522 3433 1538
rect 3454 1532 3457 1548
rect 3438 1522 3441 1528
rect 3382 1508 3393 1511
rect 3302 1492 3305 1498
rect 3306 1478 3310 1481
rect 3318 1472 3321 1488
rect 3382 1482 3385 1508
rect 3390 1482 3393 1498
rect 3422 1492 3425 1498
rect 3334 1472 3337 1478
rect 3350 1472 3353 1478
rect 3382 1472 3385 1478
rect 3410 1468 3414 1471
rect 3294 1462 3297 1468
rect 3326 1462 3329 1468
rect 3342 1462 3345 1468
rect 3358 1462 3361 1468
rect 3374 1462 3377 1468
rect 3274 1458 3278 1461
rect 3414 1452 3417 1458
rect 3422 1452 3425 1478
rect 3438 1462 3441 1488
rect 3446 1452 3449 1468
rect 3354 1448 3358 1451
rect 3390 1442 3393 1448
rect 3274 1388 3278 1391
rect 3318 1362 3321 1368
rect 3366 1362 3369 1398
rect 3382 1372 3385 1438
rect 3406 1392 3409 1438
rect 3338 1358 3342 1361
rect 3382 1352 3385 1368
rect 3394 1348 3398 1351
rect 3166 1332 3169 1338
rect 3150 1302 3153 1328
rect 3146 1288 3150 1291
rect 3094 1212 3097 1258
rect 3102 1222 3105 1258
rect 3126 1252 3129 1278
rect 3134 1272 3137 1288
rect 3174 1272 3177 1288
rect 3182 1262 3185 1268
rect 3230 1262 3233 1348
rect 3258 1338 3262 1341
rect 3238 1292 3241 1318
rect 3262 1292 3265 1298
rect 3114 1248 3118 1251
rect 3162 1248 3166 1251
rect 3126 1192 3129 1208
rect 3150 1172 3153 1248
rect 3174 1192 3177 1258
rect 3214 1242 3217 1248
rect 3230 1232 3233 1238
rect 3078 1158 3086 1161
rect 3170 1158 3174 1161
rect 3102 1152 3105 1158
rect 3134 1152 3137 1158
rect 3074 1148 3078 1151
rect 3046 1142 3049 1148
rect 3110 1142 3113 1148
rect 3078 1132 3081 1138
rect 3094 1132 3097 1138
rect 3118 1112 3121 1128
rect 3134 1102 3137 1138
rect 3142 1102 3145 1148
rect 3150 1142 3153 1158
rect 3190 1152 3193 1178
rect 3198 1152 3201 1218
rect 3238 1192 3241 1258
rect 3214 1182 3217 1188
rect 3222 1152 3225 1188
rect 3246 1182 3249 1268
rect 3254 1252 3257 1268
rect 3246 1162 3249 1178
rect 3250 1148 3254 1151
rect 3158 1122 3161 1128
rect 3094 1072 3097 1078
rect 3110 1072 3113 1078
rect 3182 1062 3185 1068
rect 3110 1012 3113 1058
rect 3142 1031 3145 1050
rect 3086 962 3089 1008
rect 3094 962 3097 988
rect 3086 952 3089 958
rect 3046 922 3049 938
rect 2946 918 2950 921
rect 2952 903 2954 907
rect 2958 903 2961 907
rect 2965 903 2968 907
rect 3054 892 3057 898
rect 2858 868 2862 871
rect 2942 862 2945 878
rect 2966 872 2969 888
rect 2978 878 2982 881
rect 3046 872 3049 888
rect 3078 872 3081 878
rect 3010 868 3014 871
rect 2870 852 2873 858
rect 2918 852 2921 858
rect 2898 848 2902 851
rect 2946 848 2950 851
rect 2806 760 2809 779
rect 2774 742 2777 748
rect 2814 741 2817 748
rect 2806 738 2817 741
rect 2838 742 2841 818
rect 2878 782 2881 818
rect 2846 752 2849 768
rect 2878 752 2881 778
rect 2894 762 2897 808
rect 2958 762 2961 858
rect 2982 762 2985 868
rect 3086 861 3089 948
rect 3094 872 3097 878
rect 3102 872 3105 908
rect 3110 892 3113 998
rect 3158 982 3161 988
rect 3118 962 3121 968
rect 3166 962 3169 968
rect 3130 948 3134 951
rect 3146 938 3150 941
rect 3126 932 3129 938
rect 3110 882 3113 888
rect 3118 882 3121 888
rect 3134 872 3137 938
rect 3142 862 3145 888
rect 3086 858 3097 861
rect 2990 852 2993 858
rect 3038 852 3041 858
rect 3070 852 3073 858
rect 3022 842 3025 848
rect 3038 802 3041 848
rect 3054 832 3057 848
rect 3082 828 3086 831
rect 3050 788 3054 791
rect 2890 758 2894 761
rect 2906 758 2921 761
rect 2918 752 2921 758
rect 2906 748 2910 751
rect 2858 738 2862 741
rect 2926 741 2929 748
rect 2922 738 2929 741
rect 2758 732 2761 738
rect 2694 652 2697 688
rect 2710 662 2713 728
rect 2718 672 2721 718
rect 2726 662 2729 708
rect 2790 672 2793 678
rect 2762 668 2766 671
rect 2794 668 2798 671
rect 2582 562 2585 588
rect 2590 562 2593 648
rect 2638 642 2641 648
rect 2610 558 2614 561
rect 2622 552 2625 618
rect 2670 562 2673 618
rect 2646 552 2649 558
rect 2478 472 2481 538
rect 2518 492 2521 528
rect 2558 482 2561 498
rect 2550 472 2553 478
rect 2538 468 2542 471
rect 2486 462 2489 468
rect 2510 462 2513 468
rect 2458 458 2462 461
rect 2440 403 2442 407
rect 2446 403 2449 407
rect 2453 403 2456 407
rect 2462 391 2465 408
rect 2454 388 2465 391
rect 2414 342 2417 348
rect 2430 342 2433 348
rect 2446 282 2449 358
rect 2454 342 2457 388
rect 2462 342 2465 378
rect 2478 372 2481 458
rect 2506 448 2510 451
rect 2518 442 2521 468
rect 2582 462 2585 548
rect 2590 462 2593 548
rect 2618 538 2622 541
rect 2666 540 2670 543
rect 2678 542 2681 558
rect 2686 542 2689 578
rect 2710 571 2713 618
rect 2734 582 2737 668
rect 2750 662 2753 668
rect 2794 658 2798 661
rect 2758 652 2761 658
rect 2750 602 2753 618
rect 2702 568 2713 571
rect 2702 562 2705 568
rect 2714 558 2718 561
rect 2730 548 2734 551
rect 2722 538 2726 541
rect 2526 452 2529 458
rect 2534 452 2537 458
rect 2570 448 2574 451
rect 2514 368 2518 371
rect 2486 352 2489 368
rect 2502 352 2505 358
rect 2474 348 2478 351
rect 2494 332 2497 338
rect 2486 312 2489 318
rect 2446 272 2449 278
rect 2494 272 2497 278
rect 2482 268 2486 271
rect 2502 262 2505 348
rect 2526 342 2529 388
rect 2534 362 2537 368
rect 2546 348 2550 351
rect 2558 342 2561 378
rect 2574 362 2577 368
rect 2582 362 2585 398
rect 2566 342 2569 348
rect 2518 338 2526 341
rect 2518 272 2521 338
rect 2526 272 2529 308
rect 2534 272 2537 298
rect 2562 278 2566 281
rect 2582 281 2585 318
rect 2574 278 2585 281
rect 2542 262 2545 268
rect 2422 258 2430 261
rect 2466 258 2470 261
rect 2514 258 2518 261
rect 2350 252 2353 258
rect 2330 248 2334 251
rect 2410 248 2414 251
rect 2262 192 2265 198
rect 2230 142 2233 148
rect 2254 92 2257 168
rect 2286 152 2289 198
rect 2398 182 2401 218
rect 2390 160 2393 179
rect 2286 92 2289 148
rect 2358 132 2361 138
rect 2342 122 2345 128
rect 2318 92 2321 108
rect 2350 92 2353 108
rect 2254 72 2257 88
rect 2382 82 2385 88
rect 2398 82 2401 148
rect 2406 92 2409 238
rect 2422 192 2425 258
rect 2478 252 2481 258
rect 2434 248 2438 251
rect 2462 222 2465 248
rect 2502 222 2505 258
rect 2514 248 2518 251
rect 2440 203 2442 207
rect 2446 203 2449 207
rect 2453 203 2456 207
rect 2422 141 2425 188
rect 2462 152 2465 198
rect 2470 142 2473 178
rect 2494 152 2497 198
rect 2502 142 2505 178
rect 2418 138 2425 141
rect 2434 138 2438 141
rect 2458 138 2462 141
rect 2414 72 2417 138
rect 2438 82 2441 138
rect 2502 132 2505 138
rect 2482 128 2486 131
rect 2526 82 2529 218
rect 2542 202 2545 218
rect 2566 182 2569 278
rect 2534 162 2537 178
rect 2554 148 2558 151
rect 2534 122 2537 148
rect 2550 138 2558 141
rect 2550 132 2553 138
rect 2566 132 2569 148
rect 2574 142 2577 278
rect 2590 272 2593 448
rect 2598 352 2601 538
rect 2626 528 2630 531
rect 2686 531 2689 538
rect 2678 528 2689 531
rect 2658 518 2662 521
rect 2606 452 2609 518
rect 2610 438 2614 441
rect 2598 342 2601 348
rect 2606 342 2609 348
rect 2622 342 2625 358
rect 2630 352 2633 518
rect 2638 412 2641 518
rect 2678 502 2681 528
rect 2698 518 2702 521
rect 2710 512 2713 518
rect 2686 482 2689 498
rect 2702 472 2705 488
rect 2646 462 2649 468
rect 2638 362 2641 388
rect 2654 352 2657 378
rect 2686 362 2689 438
rect 2702 362 2705 388
rect 2662 342 2665 348
rect 2686 342 2689 358
rect 2718 352 2721 368
rect 2698 348 2702 351
rect 2726 341 2729 408
rect 2734 352 2737 468
rect 2742 462 2745 548
rect 2750 522 2753 528
rect 2750 422 2753 448
rect 2758 362 2761 618
rect 2766 472 2769 518
rect 2774 472 2777 578
rect 2782 572 2785 648
rect 2798 642 2801 648
rect 2782 542 2785 548
rect 2790 542 2793 608
rect 2806 552 2809 738
rect 2822 662 2825 708
rect 2846 682 2849 698
rect 2830 662 2833 668
rect 2846 661 2849 678
rect 2854 672 2857 678
rect 2846 658 2854 661
rect 2838 652 2841 658
rect 2818 648 2822 651
rect 2818 558 2822 561
rect 2802 538 2806 541
rect 2822 522 2825 548
rect 2846 532 2849 658
rect 2854 542 2857 588
rect 2842 528 2846 531
rect 2794 488 2798 491
rect 2798 472 2801 478
rect 2814 471 2817 518
rect 2814 468 2825 471
rect 2770 458 2774 461
rect 2806 442 2809 468
rect 2822 462 2825 468
rect 2814 451 2817 458
rect 2838 452 2841 518
rect 2854 492 2857 538
rect 2814 448 2822 451
rect 2806 402 2809 438
rect 2766 392 2769 398
rect 2726 338 2734 341
rect 2610 328 2614 331
rect 2622 302 2625 338
rect 2638 332 2641 338
rect 2702 332 2705 338
rect 2674 328 2678 331
rect 2678 312 2681 318
rect 2602 288 2606 291
rect 2590 232 2593 258
rect 2574 132 2577 138
rect 2234 68 2238 71
rect 2322 68 2326 71
rect 2486 62 2489 78
rect 2542 72 2545 108
rect 2582 62 2585 198
rect 2610 178 2614 181
rect 2590 132 2593 178
rect 2614 132 2617 148
rect 2622 142 2625 298
rect 2686 282 2689 288
rect 2734 272 2737 338
rect 2646 202 2649 258
rect 2702 252 2705 268
rect 2742 262 2745 288
rect 2750 262 2753 318
rect 2798 312 2801 318
rect 2798 272 2801 308
rect 2806 292 2809 348
rect 2862 342 2865 718
rect 2870 692 2873 738
rect 2878 682 2881 738
rect 2910 732 2913 738
rect 2926 692 2929 728
rect 2934 682 2937 738
rect 2878 582 2881 678
rect 2914 668 2918 671
rect 2886 662 2889 668
rect 2942 662 2945 758
rect 2966 742 2969 758
rect 2982 752 2985 758
rect 2998 732 3001 748
rect 3038 742 3041 748
rect 3046 742 3049 778
rect 3094 752 3097 858
rect 3166 831 3169 918
rect 3182 892 3185 1058
rect 3190 942 3193 1138
rect 3198 1102 3201 1138
rect 3206 1132 3209 1138
rect 3198 1072 3201 1098
rect 3210 1078 3214 1081
rect 3222 1072 3225 1148
rect 3262 1142 3265 1178
rect 3230 1132 3233 1138
rect 3238 1122 3241 1128
rect 3246 1092 3249 1098
rect 3254 1082 3257 1138
rect 3202 1058 3206 1061
rect 3222 1052 3225 1058
rect 3238 1031 3241 1068
rect 3262 1062 3265 1068
rect 3270 1062 3273 1348
rect 3310 1342 3313 1348
rect 3282 1338 3286 1341
rect 3294 1332 3297 1338
rect 3334 1332 3337 1348
rect 3346 1338 3350 1341
rect 3370 1338 3374 1341
rect 3358 1332 3361 1338
rect 3294 1271 3297 1298
rect 3306 1278 3310 1281
rect 3398 1281 3401 1338
rect 3394 1278 3401 1281
rect 3294 1268 3302 1271
rect 3278 1262 3281 1268
rect 3278 1192 3281 1198
rect 3286 1182 3289 1268
rect 3318 1262 3321 1268
rect 3326 1262 3329 1278
rect 3358 1272 3361 1278
rect 3374 1272 3377 1278
rect 3382 1272 3385 1278
rect 3414 1272 3417 1298
rect 3422 1292 3425 1328
rect 3422 1272 3425 1278
rect 3350 1262 3353 1268
rect 3310 1252 3313 1258
rect 3330 1248 3334 1251
rect 3346 1248 3350 1251
rect 3286 1152 3289 1168
rect 3294 1152 3297 1188
rect 3302 1142 3305 1228
rect 3326 1152 3329 1158
rect 3278 1132 3281 1138
rect 3318 1132 3321 1148
rect 3334 1142 3337 1178
rect 3358 1152 3361 1228
rect 3366 1142 3369 1258
rect 3378 1248 3382 1251
rect 3386 1238 3390 1241
rect 3398 1212 3401 1268
rect 3406 1262 3409 1268
rect 3374 1192 3377 1198
rect 3406 1192 3409 1258
rect 3398 1188 3406 1191
rect 3350 1132 3353 1138
rect 3374 1132 3377 1148
rect 3286 1092 3289 1118
rect 3230 1028 3241 1031
rect 3197 942 3200 948
rect 3198 892 3201 918
rect 3230 902 3233 1028
rect 3270 992 3273 1058
rect 3294 1052 3297 1118
rect 3342 1082 3345 1118
rect 3350 1092 3353 1108
rect 3306 1068 3310 1071
rect 3330 1068 3334 1071
rect 3362 1068 3366 1071
rect 3338 1058 3342 1061
rect 3370 1058 3374 1061
rect 3382 1052 3385 1168
rect 3398 1132 3401 1188
rect 3418 1148 3422 1151
rect 3414 1132 3417 1138
rect 3398 1082 3401 1108
rect 3410 1068 3414 1071
rect 3430 1062 3433 1428
rect 3454 1422 3457 1478
rect 3462 1412 3465 1548
rect 3526 1532 3529 1538
rect 3514 1528 3518 1531
rect 3474 1518 3478 1521
rect 3498 1518 3502 1521
rect 3510 1472 3513 1528
rect 3534 1522 3537 1668
rect 3550 1652 3553 1668
rect 3574 1662 3577 1668
rect 3622 1662 3625 1668
rect 3618 1658 3622 1661
rect 3566 1651 3569 1658
rect 3566 1648 3574 1651
rect 3626 1648 3630 1651
rect 3606 1612 3609 1628
rect 3638 1602 3641 1668
rect 3646 1662 3649 1668
rect 3646 1582 3649 1588
rect 3578 1578 3582 1581
rect 3654 1572 3657 1668
rect 3662 1662 3665 1678
rect 3702 1672 3705 1698
rect 3734 1682 3737 1718
rect 3838 1712 3841 1848
rect 3922 1838 3926 1841
rect 3866 1818 3870 1821
rect 3926 1802 3929 1818
rect 3894 1742 3897 1798
rect 3926 1760 3929 1779
rect 3942 1752 3945 1858
rect 4014 1852 4017 1928
rect 4046 1882 4049 1918
rect 4022 1862 4025 1868
rect 4002 1848 4006 1851
rect 3950 1782 3953 1838
rect 3990 1792 3993 1838
rect 3878 1702 3881 1728
rect 3934 1712 3937 1748
rect 3830 1682 3833 1688
rect 3754 1678 3758 1681
rect 3734 1672 3737 1678
rect 3678 1652 3681 1658
rect 3694 1652 3697 1668
rect 3730 1658 3734 1661
rect 3662 1642 3665 1648
rect 3678 1612 3681 1648
rect 3710 1642 3713 1658
rect 3846 1652 3849 1668
rect 3886 1662 3889 1708
rect 3958 1662 3961 1748
rect 3930 1658 3934 1661
rect 3722 1648 3726 1651
rect 3878 1622 3881 1650
rect 3886 1612 3889 1658
rect 3946 1648 3950 1651
rect 3682 1608 3689 1611
rect 3618 1558 3622 1561
rect 3634 1558 3638 1561
rect 3554 1548 3558 1551
rect 3542 1532 3545 1548
rect 3582 1541 3585 1548
rect 3582 1538 3590 1541
rect 3558 1522 3561 1538
rect 3574 1532 3577 1538
rect 3586 1528 3590 1531
rect 3598 1522 3601 1528
rect 3534 1482 3537 1488
rect 3558 1472 3561 1478
rect 3574 1472 3577 1508
rect 3606 1492 3609 1548
rect 3630 1542 3633 1548
rect 3662 1542 3665 1568
rect 3670 1552 3673 1558
rect 3654 1532 3657 1538
rect 3654 1492 3657 1508
rect 3678 1492 3681 1598
rect 3686 1562 3689 1608
rect 3838 1592 3841 1608
rect 3694 1562 3697 1568
rect 3718 1552 3721 1578
rect 3782 1552 3785 1558
rect 3730 1548 3737 1551
rect 3734 1542 3737 1548
rect 3766 1542 3769 1548
rect 3790 1542 3793 1578
rect 3814 1552 3817 1588
rect 3918 1582 3921 1648
rect 3966 1642 3969 1778
rect 4022 1772 4025 1798
rect 4030 1792 4033 1838
rect 4062 1832 4065 1918
rect 4070 1882 4073 1928
rect 4086 1922 4089 1928
rect 4082 1878 4086 1881
rect 4094 1881 4097 1948
rect 4102 1912 4105 1948
rect 4110 1942 4113 1958
rect 4126 1952 4129 2018
rect 4134 2012 4137 2118
rect 4150 2092 4153 2098
rect 4142 2052 4145 2058
rect 4150 2042 4153 2048
rect 4138 1968 4142 1971
rect 4150 1962 4153 1978
rect 4158 1962 4161 2068
rect 4166 2062 4169 2128
rect 4190 2082 4193 2088
rect 4174 2072 4177 2078
rect 4166 1982 4169 2058
rect 4198 1962 4201 2098
rect 4206 2072 4209 2268
rect 4214 2162 4217 2178
rect 4222 2151 4225 2268
rect 4242 2258 4246 2261
rect 4230 2162 4233 2168
rect 4254 2152 4257 2268
rect 4262 2262 4265 2288
rect 4286 2272 4289 2308
rect 4310 2282 4313 2298
rect 4318 2292 4321 2348
rect 4334 2342 4337 2448
rect 4342 2442 4345 2458
rect 4366 2452 4369 2488
rect 4382 2462 4385 2538
rect 4390 2472 4393 2528
rect 4374 2372 4377 2458
rect 4382 2452 4385 2458
rect 4386 2358 4390 2361
rect 4342 2352 4345 2358
rect 4358 2342 4361 2358
rect 4370 2348 4374 2351
rect 4330 2338 4334 2341
rect 4350 2312 4353 2318
rect 4298 2278 4302 2281
rect 4290 2268 4294 2271
rect 4318 2262 4321 2288
rect 4350 2282 4353 2298
rect 4290 2258 4294 2261
rect 4270 2162 4273 2258
rect 4222 2148 4230 2151
rect 4222 2142 4225 2148
rect 4238 2142 4241 2148
rect 4246 2122 4249 2138
rect 4262 2082 4265 2158
rect 4278 2142 4281 2148
rect 4326 2142 4329 2278
rect 4338 2268 4342 2271
rect 4350 2152 4353 2218
rect 4358 2192 4361 2318
rect 4366 2272 4369 2278
rect 4374 2262 4377 2308
rect 4382 2142 4385 2338
rect 4270 2112 4273 2118
rect 4278 2092 4281 2128
rect 4298 2118 4302 2121
rect 4250 2078 4254 2081
rect 4242 2068 4246 2071
rect 4206 2052 4209 2058
rect 4262 2052 4265 2078
rect 4270 2042 4273 2058
rect 4294 2052 4297 2098
rect 4326 2082 4329 2138
rect 4358 2072 4361 2098
rect 4382 2092 4385 2128
rect 4390 2082 4393 2228
rect 4330 2068 4334 2071
rect 4318 2061 4321 2068
rect 4318 2058 4326 2061
rect 4354 2058 4358 2061
rect 4302 2052 4305 2058
rect 4230 1992 4233 1998
rect 4214 1972 4217 1978
rect 4234 1968 4238 1971
rect 4254 1962 4257 2018
rect 4278 1992 4281 2038
rect 4294 1982 4297 2048
rect 4334 2042 4337 2048
rect 4302 2032 4305 2038
rect 4270 1962 4273 1968
rect 4146 1948 4150 1951
rect 4158 1932 4161 1958
rect 4250 1948 4257 1951
rect 4166 1942 4169 1948
rect 4198 1942 4201 1948
rect 4214 1942 4217 1948
rect 4178 1938 4182 1941
rect 4222 1932 4225 1938
rect 4186 1928 4190 1931
rect 4094 1878 4102 1881
rect 4086 1862 4089 1868
rect 4074 1858 4078 1861
rect 4122 1858 4126 1861
rect 4110 1852 4113 1858
rect 4058 1818 4062 1821
rect 4038 1792 4041 1818
rect 3978 1758 3982 1761
rect 3990 1752 3993 1758
rect 3998 1712 4001 1768
rect 4038 1762 4041 1768
rect 4046 1762 4049 1798
rect 4062 1772 4065 1798
rect 3976 1703 3978 1707
rect 3982 1703 3985 1707
rect 3989 1703 3992 1707
rect 4006 1662 4009 1758
rect 4054 1752 4057 1758
rect 4022 1692 4025 1748
rect 4054 1662 4057 1718
rect 4062 1712 4065 1768
rect 4070 1682 4073 1818
rect 4098 1788 4102 1791
rect 4086 1772 4089 1788
rect 4102 1762 4105 1768
rect 4118 1762 4121 1858
rect 4142 1852 4145 1868
rect 4150 1862 4153 1888
rect 4190 1872 4193 1928
rect 4234 1878 4238 1881
rect 4246 1872 4249 1898
rect 4234 1858 4238 1861
rect 4178 1838 4182 1841
rect 4126 1802 4129 1838
rect 4126 1772 4129 1778
rect 4134 1762 4137 1768
rect 4142 1762 4145 1838
rect 4158 1802 4161 1838
rect 4166 1832 4169 1838
rect 4190 1831 4193 1858
rect 4246 1852 4249 1868
rect 4254 1862 4257 1948
rect 4278 1942 4281 1948
rect 4286 1922 4289 1958
rect 4294 1942 4297 1948
rect 4298 1928 4302 1931
rect 4278 1882 4281 1888
rect 4198 1842 4201 1848
rect 4182 1828 4193 1831
rect 4182 1792 4185 1828
rect 4190 1792 4193 1818
rect 4166 1772 4169 1778
rect 4154 1768 4158 1771
rect 4174 1762 4177 1768
rect 4190 1762 4193 1768
rect 4094 1742 4097 1748
rect 4102 1702 4105 1758
rect 4110 1722 4113 1758
rect 4158 1752 4161 1758
rect 4122 1748 4126 1751
rect 4078 1672 4081 1678
rect 4034 1658 4038 1661
rect 4074 1658 4078 1661
rect 4094 1652 4097 1668
rect 4134 1662 4137 1748
rect 4106 1658 4110 1661
rect 4026 1648 4030 1651
rect 4082 1648 4086 1651
rect 4122 1648 4126 1651
rect 3938 1638 3942 1641
rect 3862 1562 3865 1568
rect 3942 1562 3945 1618
rect 3950 1572 3953 1628
rect 3998 1622 4001 1648
rect 4006 1642 4009 1648
rect 4142 1642 4145 1738
rect 4166 1732 4169 1758
rect 4182 1752 4185 1758
rect 4190 1742 4193 1758
rect 4206 1752 4209 1788
rect 4214 1752 4217 1818
rect 4246 1792 4249 1838
rect 4266 1828 4270 1831
rect 4286 1792 4289 1908
rect 4302 1892 4305 1918
rect 4310 1912 4313 2038
rect 4338 1958 4342 1961
rect 4366 1952 4369 2068
rect 4366 1942 4369 1948
rect 4322 1938 4326 1941
rect 4346 1928 4350 1931
rect 4358 1922 4361 1938
rect 4310 1882 4313 1888
rect 4334 1872 4337 1918
rect 4322 1868 4326 1871
rect 4350 1862 4353 1918
rect 4382 1882 4385 2018
rect 4390 1932 4393 2078
rect 4366 1862 4369 1868
rect 4294 1832 4297 1858
rect 4278 1772 4281 1778
rect 4294 1762 4297 1778
rect 4302 1762 4305 1818
rect 4310 1792 4313 1858
rect 4342 1852 4345 1858
rect 4330 1848 4334 1851
rect 4318 1781 4321 1818
rect 4310 1778 4321 1781
rect 4310 1761 4313 1778
rect 4322 1768 4329 1771
rect 4310 1758 4321 1761
rect 4258 1748 4262 1751
rect 4302 1748 4310 1751
rect 4158 1722 4161 1728
rect 4166 1662 4169 1668
rect 4166 1652 4169 1658
rect 4154 1648 4158 1651
rect 4174 1642 4177 1708
rect 4182 1662 4185 1668
rect 4190 1652 4193 1728
rect 4214 1722 4217 1738
rect 4226 1728 4230 1731
rect 4226 1718 4230 1721
rect 4246 1712 4249 1718
rect 4230 1681 4233 1708
rect 4242 1688 4246 1691
rect 4230 1678 4241 1681
rect 4222 1672 4225 1678
rect 4198 1662 4201 1668
rect 4066 1638 4070 1641
rect 4114 1638 4118 1641
rect 4178 1638 4182 1641
rect 4014 1632 4017 1638
rect 4046 1632 4049 1638
rect 4038 1601 4041 1618
rect 4030 1598 4041 1601
rect 4030 1572 4033 1598
rect 4038 1582 4041 1588
rect 4046 1572 4049 1628
rect 3930 1558 3934 1561
rect 4042 1558 4046 1561
rect 3822 1552 3825 1558
rect 3686 1532 3689 1538
rect 3702 1532 3705 1538
rect 3718 1522 3721 1538
rect 3726 1522 3729 1538
rect 3774 1532 3777 1538
rect 3798 1532 3801 1538
rect 3746 1528 3750 1531
rect 3590 1472 3593 1478
rect 3606 1472 3609 1478
rect 3630 1472 3633 1488
rect 3706 1478 3710 1481
rect 3470 1462 3473 1468
rect 3510 1462 3513 1468
rect 3566 1462 3569 1468
rect 3622 1462 3625 1468
rect 3550 1452 3553 1458
rect 3442 1328 3446 1331
rect 3454 1292 3457 1298
rect 3462 1291 3465 1408
rect 3472 1403 3474 1407
rect 3478 1403 3481 1407
rect 3485 1403 3488 1407
rect 3494 1402 3497 1448
rect 3550 1432 3553 1448
rect 3526 1332 3529 1388
rect 3542 1342 3545 1368
rect 3574 1352 3577 1458
rect 3638 1452 3641 1468
rect 3694 1462 3697 1468
rect 3718 1462 3721 1508
rect 3738 1478 3742 1481
rect 3750 1462 3753 1508
rect 3798 1492 3801 1528
rect 3766 1482 3769 1488
rect 3778 1478 3782 1481
rect 3670 1452 3673 1458
rect 3582 1432 3585 1448
rect 3602 1418 3606 1421
rect 3462 1288 3473 1291
rect 3462 1272 3465 1278
rect 3470 1272 3473 1288
rect 3438 1262 3441 1268
rect 3446 1241 3449 1268
rect 3478 1262 3481 1298
rect 3502 1262 3505 1288
rect 3534 1272 3537 1288
rect 3582 1262 3585 1418
rect 3590 1362 3593 1388
rect 3638 1361 3641 1448
rect 3678 1442 3681 1448
rect 3726 1412 3729 1458
rect 3734 1422 3737 1428
rect 3630 1358 3641 1361
rect 3694 1362 3697 1368
rect 3614 1352 3617 1358
rect 3630 1342 3633 1358
rect 3702 1352 3705 1368
rect 3734 1361 3737 1418
rect 3742 1392 3745 1408
rect 3730 1358 3737 1361
rect 3750 1362 3753 1418
rect 3638 1342 3641 1348
rect 3670 1342 3673 1348
rect 3710 1342 3713 1348
rect 3650 1338 3654 1341
rect 3606 1262 3609 1338
rect 3694 1332 3697 1338
rect 3658 1328 3662 1331
rect 3670 1321 3673 1328
rect 3734 1322 3737 1338
rect 3766 1332 3769 1478
rect 3790 1472 3793 1478
rect 3798 1462 3801 1468
rect 3790 1442 3793 1458
rect 3806 1402 3809 1518
rect 3814 1492 3817 1518
rect 3830 1472 3833 1478
rect 3838 1462 3841 1518
rect 3846 1512 3849 1548
rect 3854 1522 3857 1538
rect 3886 1532 3889 1558
rect 3906 1548 3910 1551
rect 3914 1538 3918 1541
rect 3930 1538 3934 1541
rect 3902 1512 3905 1538
rect 3942 1522 3945 1548
rect 3990 1542 3993 1558
rect 4002 1538 4006 1541
rect 3846 1492 3849 1508
rect 3942 1482 3945 1488
rect 3958 1472 3961 1528
rect 3976 1503 3978 1507
rect 3982 1503 3985 1507
rect 3989 1503 3992 1507
rect 4006 1502 4009 1528
rect 4014 1502 4017 1558
rect 3898 1458 3902 1461
rect 3850 1448 3854 1451
rect 3774 1342 3777 1358
rect 3790 1352 3793 1358
rect 3658 1318 3673 1321
rect 3614 1292 3617 1318
rect 3726 1292 3729 1318
rect 3686 1282 3689 1288
rect 3650 1278 3654 1281
rect 3614 1272 3617 1278
rect 3694 1272 3697 1278
rect 3622 1262 3625 1268
rect 3670 1262 3673 1268
rect 3694 1262 3697 1268
rect 3702 1262 3705 1288
rect 3518 1252 3521 1258
rect 3438 1238 3449 1241
rect 3438 1192 3441 1238
rect 3498 1228 3502 1231
rect 3472 1203 3474 1207
rect 3478 1203 3481 1207
rect 3485 1203 3488 1207
rect 3510 1192 3513 1248
rect 3526 1232 3529 1258
rect 3542 1252 3545 1258
rect 3582 1252 3585 1258
rect 3606 1242 3609 1258
rect 3726 1242 3729 1278
rect 3742 1272 3745 1288
rect 3750 1272 3753 1328
rect 3758 1292 3761 1318
rect 3766 1281 3769 1328
rect 3766 1278 3774 1281
rect 3782 1272 3785 1278
rect 3790 1272 3793 1318
rect 3798 1292 3801 1358
rect 3806 1352 3809 1358
rect 3814 1341 3817 1418
rect 3822 1352 3825 1448
rect 3858 1418 3862 1421
rect 3902 1372 3905 1398
rect 3910 1392 3913 1408
rect 3934 1372 3937 1398
rect 3942 1392 3945 1438
rect 3990 1422 3993 1450
rect 4022 1412 4025 1548
rect 4054 1522 4057 1548
rect 3834 1368 3838 1371
rect 3830 1352 3833 1358
rect 3870 1342 3873 1348
rect 3878 1342 3881 1348
rect 3814 1338 3822 1341
rect 3806 1292 3809 1298
rect 3814 1282 3817 1288
rect 3822 1282 3825 1338
rect 3858 1328 3865 1331
rect 3862 1292 3865 1328
rect 3878 1282 3881 1288
rect 3826 1268 3830 1271
rect 3758 1262 3761 1268
rect 3790 1262 3793 1268
rect 3886 1262 3889 1358
rect 3894 1292 3897 1348
rect 3918 1332 3921 1358
rect 3934 1352 3937 1368
rect 3950 1362 3953 1378
rect 3958 1352 3961 1378
rect 3970 1368 3974 1371
rect 4026 1358 4030 1361
rect 4038 1352 4041 1378
rect 4046 1372 4049 1508
rect 4054 1462 4057 1518
rect 4062 1512 4065 1568
rect 4102 1562 4105 1618
rect 4118 1572 4121 1578
rect 4134 1571 4137 1618
rect 4198 1592 4201 1638
rect 4214 1622 4217 1628
rect 4222 1592 4225 1658
rect 4126 1568 4137 1571
rect 4146 1568 4150 1571
rect 4194 1568 4198 1571
rect 4086 1542 4089 1558
rect 4106 1538 4110 1541
rect 4106 1528 4113 1531
rect 4062 1472 4065 1478
rect 4062 1442 4065 1458
rect 4070 1452 4073 1498
rect 4102 1462 4105 1468
rect 4086 1452 4089 1458
rect 4110 1452 4113 1528
rect 4118 1462 4121 1468
rect 4078 1442 4081 1448
rect 4054 1392 4057 1438
rect 4086 1392 4089 1428
rect 4046 1362 4049 1368
rect 4062 1362 4065 1368
rect 4070 1352 4073 1378
rect 3994 1348 3998 1351
rect 3894 1262 3897 1268
rect 3834 1258 3838 1261
rect 3438 1182 3441 1188
rect 3510 1182 3513 1188
rect 3454 1152 3457 1178
rect 3526 1162 3529 1228
rect 3566 1192 3569 1218
rect 3590 1202 3593 1218
rect 3438 1072 3441 1078
rect 3446 1062 3449 1068
rect 3370 1048 3374 1051
rect 3286 1012 3289 1048
rect 3294 972 3297 1048
rect 3350 1042 3353 1048
rect 3326 960 3329 979
rect 3382 962 3385 1048
rect 3390 1012 3393 1018
rect 3238 952 3241 958
rect 3294 942 3297 948
rect 3398 942 3401 948
rect 3366 932 3369 938
rect 3222 872 3225 878
rect 3246 872 3249 878
rect 3174 842 3177 858
rect 3166 828 3174 831
rect 3134 772 3137 818
rect 3166 802 3169 818
rect 3182 760 3185 779
rect 3190 761 3193 868
rect 3190 758 3198 761
rect 3010 738 3014 741
rect 3014 722 3017 728
rect 3094 722 3097 748
rect 3150 742 3153 748
rect 2986 718 2990 721
rect 2952 703 2954 707
rect 2958 703 2961 707
rect 2965 703 2968 707
rect 2958 662 2961 678
rect 2966 672 2969 688
rect 2974 672 2977 718
rect 3022 692 3025 718
rect 3026 678 3030 681
rect 3010 668 3014 671
rect 3070 662 3073 718
rect 3134 712 3137 728
rect 3002 658 3006 661
rect 3066 658 3070 661
rect 2910 632 2913 658
rect 2950 652 2953 658
rect 2986 648 2990 651
rect 3006 642 3009 648
rect 2890 588 2894 591
rect 3022 560 3025 579
rect 3038 552 3041 658
rect 3110 632 3113 678
rect 3126 672 3129 698
rect 3198 682 3201 758
rect 3206 692 3209 868
rect 3242 858 3246 861
rect 3214 832 3217 858
rect 3226 848 3230 851
rect 3222 752 3225 798
rect 3254 792 3257 868
rect 3262 862 3265 908
rect 3278 902 3281 928
rect 3286 862 3289 908
rect 3310 882 3313 888
rect 3262 852 3265 858
rect 3278 842 3281 848
rect 3246 742 3249 788
rect 3270 742 3273 758
rect 3294 752 3297 768
rect 3310 752 3313 818
rect 3318 812 3321 848
rect 3326 792 3329 928
rect 3374 882 3377 918
rect 3382 882 3385 908
rect 3342 872 3345 878
rect 3390 871 3393 918
rect 3406 912 3409 948
rect 3422 942 3425 948
rect 3414 932 3417 938
rect 3390 868 3398 871
rect 3334 862 3337 868
rect 3342 851 3345 858
rect 3338 848 3345 851
rect 3350 782 3353 868
rect 3390 862 3393 868
rect 3414 862 3417 908
rect 3430 882 3433 1058
rect 3438 952 3441 978
rect 3454 972 3457 1148
rect 3478 1142 3481 1158
rect 3494 1142 3497 1148
rect 3466 1128 3470 1131
rect 3502 1131 3505 1138
rect 3494 1128 3505 1131
rect 3462 1092 3465 1108
rect 3474 1078 3478 1081
rect 3466 1048 3470 1051
rect 3482 1048 3486 1051
rect 3494 1032 3497 1128
rect 3522 1118 3526 1121
rect 3510 1072 3513 1078
rect 3518 1072 3521 1088
rect 3534 1062 3537 1158
rect 3622 1152 3625 1218
rect 3654 1192 3657 1218
rect 3670 1202 3673 1218
rect 3670 1162 3673 1188
rect 3702 1182 3705 1218
rect 3726 1162 3729 1238
rect 3750 1202 3753 1258
rect 3846 1252 3849 1258
rect 3902 1252 3905 1308
rect 3926 1292 3929 1348
rect 3910 1262 3913 1288
rect 3922 1278 3926 1281
rect 3942 1262 3945 1288
rect 3922 1238 3926 1241
rect 3934 1232 3937 1248
rect 3950 1242 3953 1348
rect 3966 1292 3969 1348
rect 4022 1342 4025 1348
rect 4026 1328 4030 1331
rect 3976 1303 3978 1307
rect 3982 1303 3985 1307
rect 3989 1303 3992 1307
rect 3998 1262 4001 1268
rect 4006 1252 4009 1328
rect 4022 1272 4025 1278
rect 4050 1258 4054 1261
rect 4014 1252 4017 1258
rect 4022 1252 4025 1258
rect 4042 1248 4046 1251
rect 3766 1172 3769 1218
rect 3806 1162 3809 1178
rect 3706 1158 3710 1161
rect 3674 1148 3678 1151
rect 3722 1148 3726 1151
rect 3746 1148 3750 1151
rect 3606 1132 3609 1148
rect 3622 1112 3625 1138
rect 3698 1128 3702 1131
rect 3550 1071 3553 1098
rect 3558 1092 3561 1108
rect 3578 1078 3582 1081
rect 3626 1078 3630 1081
rect 3566 1072 3569 1078
rect 3654 1072 3657 1098
rect 3694 1082 3697 1118
rect 3710 1112 3713 1118
rect 3718 1092 3721 1128
rect 3702 1082 3705 1088
rect 3666 1078 3670 1081
rect 3726 1072 3729 1108
rect 3734 1092 3737 1138
rect 3758 1132 3761 1158
rect 3822 1152 3825 1208
rect 3862 1162 3865 1218
rect 3846 1152 3849 1158
rect 3778 1148 3782 1151
rect 3798 1142 3801 1148
rect 3770 1138 3774 1141
rect 3826 1138 3830 1141
rect 3742 1102 3745 1128
rect 3766 1092 3769 1118
rect 3790 1082 3793 1138
rect 3814 1132 3817 1138
rect 3838 1132 3841 1138
rect 3886 1132 3889 1138
rect 3862 1128 3870 1131
rect 3862 1122 3865 1128
rect 3882 1118 3886 1121
rect 3838 1082 3841 1088
rect 3550 1068 3558 1071
rect 3626 1068 3630 1071
rect 3658 1068 3662 1071
rect 3722 1068 3726 1071
rect 3738 1068 3742 1071
rect 3542 1062 3545 1068
rect 3598 1062 3601 1068
rect 3646 1062 3649 1068
rect 3686 1062 3689 1068
rect 3506 1058 3510 1061
rect 3570 1058 3574 1061
rect 3666 1058 3670 1061
rect 3794 1058 3798 1061
rect 3472 1003 3474 1007
rect 3478 1003 3481 1007
rect 3485 1003 3488 1007
rect 3494 962 3497 1028
rect 3502 952 3505 1048
rect 3526 972 3529 1018
rect 3534 992 3537 1058
rect 3542 992 3545 1058
rect 3602 1048 3606 1051
rect 3558 992 3561 1038
rect 3510 952 3513 958
rect 3518 952 3521 968
rect 3474 948 3478 951
rect 3462 942 3465 948
rect 3450 938 3454 941
rect 3438 892 3441 938
rect 3518 932 3521 938
rect 3458 928 3462 931
rect 3438 882 3441 888
rect 3422 872 3425 878
rect 3434 868 3438 871
rect 3446 862 3449 918
rect 3526 872 3529 968
rect 3558 942 3561 988
rect 3574 962 3577 1008
rect 3662 992 3665 1028
rect 3594 958 3598 961
rect 3546 938 3550 941
rect 3538 888 3542 891
rect 3466 868 3470 871
rect 3362 858 3366 861
rect 3402 858 3406 861
rect 3358 832 3361 838
rect 3278 742 3281 748
rect 3286 742 3289 748
rect 3422 742 3425 828
rect 3454 762 3457 868
rect 3478 862 3481 868
rect 3506 858 3510 861
rect 3518 852 3521 858
rect 3502 842 3505 848
rect 3470 832 3473 838
rect 3472 803 3474 807
rect 3478 803 3481 807
rect 3485 803 3488 807
rect 3470 762 3473 788
rect 3494 762 3497 798
rect 3298 738 3302 741
rect 3222 732 3225 738
rect 3174 622 3177 648
rect 3198 592 3201 678
rect 3214 652 3217 668
rect 3230 662 3233 698
rect 3238 692 3241 728
rect 3310 722 3313 728
rect 3302 682 3305 718
rect 3334 682 3337 698
rect 3406 692 3409 728
rect 3422 711 3425 718
rect 3414 708 3425 711
rect 3342 682 3345 688
rect 3358 682 3361 688
rect 3250 678 3254 681
rect 3222 642 3225 658
rect 3254 652 3257 658
rect 2930 548 2934 551
rect 2990 542 2993 548
rect 3062 542 3065 588
rect 3070 582 3073 588
rect 3086 542 3089 588
rect 3110 568 3126 571
rect 3110 552 3113 568
rect 3126 552 3129 558
rect 3094 542 3097 548
rect 3118 542 3121 548
rect 2974 532 2977 538
rect 2878 482 2881 518
rect 2952 503 2954 507
rect 2958 503 2961 507
rect 2965 503 2968 507
rect 2934 482 2937 498
rect 2934 472 2937 478
rect 2950 472 2953 488
rect 2894 352 2897 458
rect 2982 431 2985 450
rect 2910 362 2913 388
rect 2978 358 2982 361
rect 3002 358 3006 361
rect 3014 352 3017 508
rect 3070 482 3073 518
rect 3110 492 3113 538
rect 3106 478 3110 481
rect 3062 472 3065 478
rect 3094 472 3097 478
rect 3042 468 3046 471
rect 3122 468 3126 471
rect 3134 462 3137 548
rect 3150 532 3153 548
rect 3166 542 3169 558
rect 3174 552 3177 578
rect 3190 552 3193 558
rect 3178 538 3182 541
rect 3206 532 3209 558
rect 3222 552 3225 638
rect 3230 612 3233 618
rect 3254 572 3257 618
rect 3214 542 3217 548
rect 3230 541 3233 558
rect 3226 538 3233 541
rect 3238 532 3241 538
rect 3230 522 3233 528
rect 3206 482 3209 518
rect 3246 512 3249 548
rect 3254 542 3257 548
rect 3270 542 3273 678
rect 3298 668 3302 671
rect 3330 668 3334 671
rect 3362 658 3366 661
rect 3386 658 3390 661
rect 3398 661 3401 688
rect 3414 672 3417 708
rect 3422 672 3425 698
rect 3398 658 3406 661
rect 3386 648 3390 651
rect 3410 648 3414 651
rect 3454 642 3457 758
rect 3462 752 3465 758
rect 3510 742 3513 778
rect 3522 768 3526 771
rect 3518 752 3521 758
rect 3510 681 3513 738
rect 3510 678 3521 681
rect 3510 662 3513 668
rect 3474 658 3478 661
rect 3498 658 3502 661
rect 3494 642 3497 648
rect 3278 562 3281 618
rect 3254 491 3257 538
rect 3246 488 3257 491
rect 3162 478 3166 481
rect 3210 468 3214 471
rect 3234 468 3238 471
rect 3142 462 3145 468
rect 3166 462 3169 468
rect 3050 458 3054 461
rect 3074 458 3078 461
rect 3094 452 3097 458
rect 3158 452 3161 458
rect 3034 448 3038 451
rect 3046 352 3049 418
rect 3062 352 3065 358
rect 2846 311 2849 328
rect 2846 308 2857 311
rect 2814 292 2817 298
rect 2806 272 2809 278
rect 2846 272 2849 298
rect 2790 262 2793 268
rect 2774 252 2777 258
rect 2750 222 2753 248
rect 2630 152 2633 178
rect 2662 152 2665 178
rect 2718 172 2721 198
rect 2650 138 2654 141
rect 2590 122 2593 128
rect 2590 82 2593 118
rect 2622 92 2625 138
rect 2638 132 2641 138
rect 2678 122 2681 128
rect 2638 112 2641 118
rect 2610 78 2614 81
rect 2614 72 2617 78
rect 2630 72 2633 78
rect 2662 62 2665 78
rect 2670 72 2673 88
rect 2678 72 2681 78
rect 2678 62 2681 68
rect 2686 62 2689 158
rect 2702 152 2705 158
rect 2718 152 2721 168
rect 2694 72 2697 148
rect 2726 142 2729 178
rect 2750 162 2753 208
rect 2774 142 2777 148
rect 2782 142 2785 258
rect 2822 242 2825 248
rect 2806 162 2809 188
rect 2738 138 2742 141
rect 2702 92 2705 98
rect 1562 58 1566 61
rect 1770 58 1774 61
rect 1834 58 1838 61
rect 2002 58 2006 61
rect 2218 58 2222 61
rect 2274 58 2278 61
rect 2306 58 2310 61
rect 2338 58 2342 61
rect 2362 58 2366 61
rect 2650 58 2654 61
rect 1470 31 1473 50
rect 1598 -18 1601 48
rect 1750 31 1753 50
rect 2010 48 2014 51
rect 1942 22 1945 48
rect 2038 42 2041 48
rect 2022 -18 2025 38
rect 2134 12 2137 48
rect 2154 38 2158 41
rect 2174 31 2177 48
rect 2170 28 2177 31
rect 2134 -18 2137 8
rect 2150 -18 2153 8
rect 2166 -18 2169 28
rect 2270 -18 2273 58
rect 2622 52 2625 58
rect 2702 52 2705 88
rect 2734 82 2737 138
rect 2766 132 2769 138
rect 2774 72 2777 138
rect 2790 92 2793 98
rect 2710 62 2713 68
rect 2758 62 2761 68
rect 2782 62 2785 78
rect 2814 62 2817 218
rect 2830 212 2833 258
rect 2838 202 2841 258
rect 2854 222 2857 308
rect 2902 262 2905 348
rect 2974 342 2977 348
rect 2962 338 2966 341
rect 2934 302 2937 318
rect 2942 312 2945 328
rect 2952 303 2954 307
rect 2958 303 2961 307
rect 2965 303 2968 307
rect 2942 282 2945 288
rect 2958 272 2961 288
rect 2866 248 2870 251
rect 2950 192 2953 208
rect 2854 132 2857 138
rect 2870 132 2873 168
rect 2910 142 2913 148
rect 2958 142 2961 258
rect 2990 222 2993 250
rect 2990 192 2993 208
rect 2998 192 3001 348
rect 3014 342 3017 348
rect 3010 338 3014 341
rect 3042 338 3046 341
rect 3022 302 3025 338
rect 3030 292 3033 318
rect 3054 302 3057 338
rect 3070 292 3073 448
rect 3090 388 3094 391
rect 3078 362 3081 378
rect 3082 338 3086 341
rect 3078 272 3081 298
rect 3066 268 3070 271
rect 3050 258 3054 261
rect 3082 258 3086 261
rect 3046 242 3049 248
rect 3062 242 3065 258
rect 3094 252 3097 258
rect 3102 252 3105 378
rect 3110 272 3113 408
rect 3174 382 3177 468
rect 3182 462 3185 468
rect 3190 452 3193 468
rect 3246 462 3249 488
rect 3234 458 3238 461
rect 3198 452 3201 458
rect 3262 452 3265 518
rect 3286 462 3289 588
rect 3310 581 3313 618
rect 3350 602 3353 618
rect 3374 612 3377 618
rect 3430 612 3433 618
rect 3472 603 3474 607
rect 3478 603 3481 607
rect 3485 603 3488 607
rect 3338 588 3342 591
rect 3302 578 3313 581
rect 3302 552 3305 578
rect 3310 552 3313 568
rect 3330 558 3334 561
rect 3438 542 3441 588
rect 3486 562 3489 588
rect 3470 552 3473 558
rect 3518 542 3521 678
rect 3534 662 3537 728
rect 3542 682 3545 728
rect 3550 672 3553 928
rect 3558 742 3561 758
rect 3566 752 3569 758
rect 3574 742 3577 958
rect 3586 948 3590 951
rect 3582 852 3585 938
rect 3606 922 3609 958
rect 3614 952 3617 978
rect 3650 948 3654 951
rect 3622 942 3625 948
rect 3638 922 3641 928
rect 3626 918 3630 921
rect 3646 901 3649 908
rect 3638 898 3649 901
rect 3622 882 3625 888
rect 3638 872 3641 898
rect 3582 782 3585 848
rect 3638 821 3641 858
rect 3638 818 3649 821
rect 3646 802 3649 818
rect 3646 792 3649 798
rect 3590 762 3593 768
rect 3598 742 3601 758
rect 3614 752 3617 768
rect 3634 748 3638 751
rect 3626 738 3630 741
rect 3558 732 3561 738
rect 3586 728 3590 731
rect 3590 682 3593 688
rect 3542 652 3545 668
rect 3550 662 3553 668
rect 3530 648 3534 651
rect 3310 532 3313 538
rect 3422 522 3425 528
rect 3302 492 3305 508
rect 3306 468 3310 471
rect 3274 458 3278 461
rect 3250 418 3254 421
rect 3214 402 3217 418
rect 3190 342 3193 388
rect 3222 360 3225 379
rect 3270 362 3273 448
rect 3274 358 3278 361
rect 3298 358 3305 361
rect 3302 352 3305 358
rect 3290 348 3294 351
rect 3118 272 3121 298
rect 3154 288 3158 291
rect 3110 262 3113 268
rect 3134 262 3137 268
rect 3142 262 3145 278
rect 3158 272 3161 288
rect 3062 162 3065 238
rect 3110 192 3113 218
rect 3126 152 3129 258
rect 3134 192 3137 248
rect 3054 142 3057 148
rect 2870 82 2873 118
rect 2886 72 2889 78
rect 2934 62 2937 138
rect 2952 103 2954 107
rect 2958 103 2961 107
rect 2965 103 2968 107
rect 3078 82 3081 88
rect 3002 78 3006 81
rect 2990 72 2993 78
rect 3094 72 3097 78
rect 2970 68 2974 71
rect 3038 62 3041 68
rect 3142 62 3145 128
rect 3174 122 3177 328
rect 3238 322 3241 348
rect 3258 338 3262 341
rect 3274 338 3278 341
rect 3298 338 3302 341
rect 3238 252 3241 278
rect 3254 272 3257 288
rect 3302 282 3305 318
rect 3310 302 3313 338
rect 3318 322 3321 518
rect 3406 482 3409 488
rect 3422 472 3425 488
rect 3510 462 3513 528
rect 3526 481 3529 648
rect 3550 612 3553 658
rect 3558 632 3561 678
rect 3566 652 3569 668
rect 3574 632 3577 658
rect 3534 552 3537 568
rect 3558 532 3561 628
rect 3566 592 3569 618
rect 3598 592 3601 718
rect 3614 671 3617 728
rect 3606 668 3617 671
rect 3630 672 3633 678
rect 3606 662 3609 668
rect 3574 542 3577 568
rect 3590 562 3593 578
rect 3582 522 3585 548
rect 3550 501 3553 518
rect 3582 512 3585 518
rect 3542 498 3553 501
rect 3526 478 3534 481
rect 3518 462 3521 468
rect 3542 462 3545 498
rect 3554 488 3558 491
rect 3334 362 3337 378
rect 3374 352 3377 358
rect 3330 348 3334 351
rect 3386 348 3390 351
rect 3342 342 3345 348
rect 3366 342 3369 348
rect 3334 292 3337 308
rect 3350 302 3353 338
rect 3302 262 3305 278
rect 3322 268 3326 271
rect 3286 231 3289 250
rect 3210 188 3214 191
rect 3186 138 3190 141
rect 3174 112 3177 118
rect 3198 72 3201 178
rect 3214 82 3217 88
rect 3222 72 3225 78
rect 3238 72 3241 228
rect 3334 152 3337 278
rect 3346 258 3350 261
rect 3350 162 3353 188
rect 3246 132 3249 148
rect 3302 142 3305 148
rect 3358 142 3361 318
rect 3382 292 3385 298
rect 3370 258 3374 261
rect 3286 132 3289 138
rect 3286 91 3289 128
rect 3366 102 3369 248
rect 3374 142 3377 158
rect 3390 152 3393 318
rect 3398 282 3401 318
rect 3414 292 3417 378
rect 3422 342 3425 458
rect 3470 422 3473 448
rect 3566 442 3569 468
rect 3574 462 3577 508
rect 3598 471 3601 518
rect 3594 468 3601 471
rect 3472 403 3474 407
rect 3478 403 3481 407
rect 3485 403 3488 407
rect 3434 388 3438 391
rect 3474 348 3478 351
rect 3414 282 3417 288
rect 3398 142 3401 268
rect 3406 262 3409 278
rect 3438 262 3441 288
rect 3478 252 3481 348
rect 3534 342 3537 398
rect 3566 360 3569 379
rect 3518 322 3521 328
rect 3486 262 3489 308
rect 3582 302 3585 468
rect 3594 458 3598 461
rect 3606 452 3609 658
rect 3614 652 3617 658
rect 3654 652 3657 778
rect 3662 752 3665 768
rect 3670 662 3673 938
rect 3678 862 3681 1058
rect 3706 1048 3710 1051
rect 3702 952 3705 1038
rect 3734 992 3737 1018
rect 3854 1002 3857 1068
rect 3886 1031 3889 1050
rect 3822 992 3825 998
rect 3718 952 3721 988
rect 3786 958 3790 961
rect 3690 918 3694 921
rect 3686 822 3689 848
rect 3690 758 3694 761
rect 3702 732 3705 948
rect 3734 942 3737 958
rect 3798 952 3801 988
rect 3850 968 3854 971
rect 3762 948 3766 951
rect 3834 948 3838 951
rect 3774 942 3777 948
rect 3746 938 3750 941
rect 3818 938 3822 941
rect 3710 932 3713 938
rect 3710 862 3713 918
rect 3726 882 3729 888
rect 3734 882 3737 938
rect 3742 922 3745 928
rect 3758 922 3761 938
rect 3806 932 3809 938
rect 3786 918 3790 921
rect 3742 902 3745 918
rect 3718 872 3721 878
rect 3738 868 3742 871
rect 3750 851 3753 918
rect 3758 862 3761 918
rect 3790 892 3793 908
rect 3782 872 3785 878
rect 3798 872 3801 888
rect 3814 872 3817 928
rect 3846 882 3849 898
rect 3810 868 3814 871
rect 3746 848 3753 851
rect 3766 852 3769 868
rect 3822 862 3825 878
rect 3862 872 3865 878
rect 3870 862 3873 968
rect 3778 858 3782 861
rect 3810 858 3814 861
rect 3834 858 3838 861
rect 3870 852 3873 858
rect 3878 852 3881 958
rect 3894 872 3897 1218
rect 3950 1162 3953 1218
rect 3990 1192 3993 1238
rect 3998 1182 4001 1218
rect 4030 1212 4033 1238
rect 4062 1212 4065 1238
rect 4078 1212 4081 1368
rect 4094 1362 4097 1438
rect 4102 1392 4105 1438
rect 4098 1348 4102 1351
rect 4094 1292 4097 1338
rect 4110 1332 4113 1448
rect 4126 1442 4129 1568
rect 4138 1558 4142 1561
rect 4142 1462 4145 1468
rect 4150 1442 4153 1548
rect 4158 1532 4161 1538
rect 4166 1522 4169 1558
rect 4174 1542 4177 1558
rect 4206 1552 4209 1558
rect 4182 1542 4185 1548
rect 4214 1542 4217 1548
rect 4162 1478 4166 1481
rect 4194 1468 4198 1471
rect 4166 1462 4169 1468
rect 4170 1448 4174 1451
rect 4182 1432 4185 1458
rect 4206 1452 4209 1488
rect 4214 1482 4217 1538
rect 4214 1462 4217 1478
rect 4222 1442 4225 1568
rect 4238 1562 4241 1678
rect 4246 1662 4249 1678
rect 4246 1562 4249 1658
rect 4254 1652 4257 1678
rect 4262 1652 4265 1658
rect 4270 1642 4273 1678
rect 4262 1601 4265 1618
rect 4254 1598 4265 1601
rect 4254 1572 4257 1598
rect 4278 1592 4281 1748
rect 4286 1652 4289 1658
rect 4294 1652 4297 1658
rect 4294 1632 4297 1638
rect 4262 1582 4265 1588
rect 4270 1562 4273 1578
rect 4294 1571 4297 1618
rect 4290 1568 4297 1571
rect 4230 1542 4233 1548
rect 4238 1502 4241 1558
rect 4274 1548 4278 1551
rect 4246 1542 4249 1548
rect 4242 1468 4246 1471
rect 4194 1438 4198 1441
rect 4214 1432 4217 1438
rect 4222 1432 4225 1438
rect 4222 1402 4225 1428
rect 4186 1388 4190 1391
rect 4126 1362 4129 1368
rect 4118 1352 4121 1358
rect 4134 1352 4137 1378
rect 4146 1368 4150 1371
rect 4154 1358 4158 1361
rect 4166 1352 4169 1378
rect 4178 1368 4182 1371
rect 4214 1362 4217 1368
rect 4190 1332 4193 1338
rect 4102 1282 4105 1298
rect 4086 1272 4089 1278
rect 4110 1242 4113 1258
rect 4110 1192 4113 1218
rect 4026 1188 4030 1191
rect 3970 1168 3974 1171
rect 4018 1168 4022 1171
rect 4050 1168 4054 1171
rect 3902 1132 3905 1158
rect 3926 1142 3929 1148
rect 3958 1142 3961 1148
rect 3902 942 3905 1078
rect 3934 1062 3937 1138
rect 3942 1112 3945 1128
rect 3946 1068 3950 1071
rect 3966 1062 3969 1168
rect 3994 1158 3998 1161
rect 4058 1158 4062 1161
rect 4030 1152 4033 1158
rect 4066 1148 4070 1151
rect 4006 1142 4009 1148
rect 4038 1142 4041 1148
rect 4086 1142 4089 1148
rect 4070 1132 4073 1138
rect 4090 1128 4094 1131
rect 4102 1121 4105 1168
rect 4118 1162 4121 1298
rect 4126 1252 4129 1328
rect 4198 1321 4201 1348
rect 4214 1342 4217 1348
rect 4190 1318 4201 1321
rect 4150 1262 4153 1318
rect 4130 1248 4134 1251
rect 4138 1248 4142 1251
rect 4162 1238 4169 1241
rect 4134 1192 4137 1228
rect 4166 1192 4169 1238
rect 4174 1222 4177 1258
rect 4182 1192 4185 1308
rect 4190 1292 4193 1318
rect 4198 1202 4201 1278
rect 4206 1252 4209 1338
rect 4214 1262 4217 1268
rect 4222 1242 4225 1398
rect 4238 1392 4241 1458
rect 4262 1422 4265 1478
rect 4278 1462 4281 1468
rect 4286 1452 4289 1518
rect 4294 1492 4297 1548
rect 4290 1448 4294 1451
rect 4230 1372 4233 1388
rect 4286 1372 4289 1448
rect 4302 1392 4305 1748
rect 4318 1702 4321 1758
rect 4318 1682 4321 1698
rect 4310 1678 4318 1681
rect 4310 1612 4313 1678
rect 4318 1662 4321 1668
rect 4326 1651 4329 1768
rect 4342 1762 4345 1768
rect 4358 1752 4361 1858
rect 4358 1692 4361 1748
rect 4350 1672 4353 1688
rect 4318 1648 4329 1651
rect 4318 1592 4321 1648
rect 4334 1642 4337 1668
rect 4342 1652 4345 1658
rect 4314 1568 4318 1571
rect 4326 1562 4329 1578
rect 4334 1562 4337 1608
rect 4342 1592 4345 1628
rect 4350 1622 4353 1658
rect 4358 1652 4361 1658
rect 4314 1548 4318 1551
rect 4342 1532 4345 1548
rect 4310 1482 4313 1488
rect 4282 1358 4286 1361
rect 4238 1312 4241 1348
rect 4246 1312 4249 1358
rect 4294 1351 4297 1368
rect 4310 1362 4313 1468
rect 4322 1458 4326 1461
rect 4342 1432 4345 1438
rect 4350 1422 4353 1568
rect 4358 1462 4361 1618
rect 4326 1392 4329 1418
rect 4338 1358 4342 1361
rect 4282 1348 4297 1351
rect 4310 1348 4318 1351
rect 4346 1348 4350 1351
rect 4254 1322 4257 1338
rect 4262 1322 4265 1348
rect 4302 1342 4305 1348
rect 4254 1272 4257 1278
rect 4230 1262 4233 1268
rect 4262 1262 4265 1308
rect 4286 1292 4289 1318
rect 4310 1292 4313 1348
rect 4358 1342 4361 1458
rect 4318 1332 4321 1338
rect 4290 1278 4294 1281
rect 4310 1268 4318 1271
rect 4270 1262 4273 1268
rect 4250 1258 4254 1261
rect 4262 1252 4265 1258
rect 4278 1251 4281 1268
rect 4270 1248 4281 1251
rect 4178 1168 4182 1171
rect 4190 1162 4193 1198
rect 4238 1192 4241 1208
rect 4246 1192 4249 1238
rect 4270 1192 4273 1248
rect 4310 1192 4313 1268
rect 4334 1262 4337 1278
rect 4326 1252 4329 1258
rect 4334 1252 4337 1258
rect 4342 1242 4345 1258
rect 4350 1242 4353 1268
rect 4366 1262 4369 1748
rect 4382 1741 4385 1828
rect 4390 1752 4393 1758
rect 4382 1738 4393 1741
rect 4374 1682 4377 1718
rect 4374 1652 4377 1658
rect 4374 1452 4377 1648
rect 4390 1462 4393 1738
rect 4374 1382 4377 1418
rect 4374 1282 4377 1338
rect 4390 1312 4393 1458
rect 4358 1252 4361 1258
rect 4214 1182 4217 1188
rect 4238 1172 4241 1188
rect 4262 1172 4265 1178
rect 4302 1172 4305 1178
rect 4326 1172 4329 1178
rect 4210 1168 4214 1171
rect 4338 1168 4342 1171
rect 4350 1162 4353 1198
rect 4358 1192 4361 1238
rect 4366 1182 4369 1258
rect 4382 1192 4385 1218
rect 4370 1168 4377 1171
rect 4218 1158 4222 1161
rect 4298 1158 4305 1161
rect 4314 1158 4318 1161
rect 4110 1152 4113 1158
rect 4150 1152 4153 1158
rect 4130 1148 4134 1151
rect 4094 1118 4105 1121
rect 4118 1138 4126 1141
rect 3976 1103 3978 1107
rect 3982 1103 3985 1107
rect 3989 1103 3992 1107
rect 4094 1092 4097 1118
rect 4118 1092 4121 1138
rect 4158 1122 4161 1158
rect 4234 1148 4241 1151
rect 4166 1142 4169 1148
rect 4198 1142 4201 1148
rect 3974 1072 3977 1078
rect 3926 972 3929 1048
rect 3942 1042 3945 1058
rect 3966 1042 3969 1048
rect 3974 1042 3977 1058
rect 3982 1052 3985 1088
rect 4130 1078 4134 1081
rect 4150 1072 4153 1078
rect 4174 1072 4177 1088
rect 4190 1082 4193 1128
rect 4198 1082 4201 1098
rect 4206 1082 4209 1088
rect 4190 1072 4193 1078
rect 4106 1068 4110 1071
rect 4166 1062 4169 1068
rect 4098 1058 4102 1061
rect 4146 1058 4150 1061
rect 4186 1058 4190 1061
rect 4014 1052 4017 1058
rect 4046 1052 4049 1058
rect 4078 1052 4081 1058
rect 4158 1052 4161 1058
rect 4198 1052 4201 1078
rect 4238 1062 4241 1148
rect 4270 1132 4273 1148
rect 4254 1092 4257 1098
rect 4262 1092 4265 1108
rect 4294 1102 4297 1148
rect 4302 1092 4305 1158
rect 4330 1148 4334 1151
rect 4326 1142 4329 1148
rect 4302 1082 4305 1088
rect 4274 1058 4278 1061
rect 3966 952 3969 988
rect 3930 948 3934 951
rect 3918 942 3921 948
rect 3954 938 3958 941
rect 3910 932 3913 938
rect 3918 892 3921 938
rect 3942 922 3945 928
rect 3982 922 3985 1048
rect 3998 992 4001 1038
rect 4006 1032 4009 1048
rect 4026 1038 4030 1041
rect 4038 1012 4041 1048
rect 4058 1038 4062 1041
rect 4070 1022 4073 1048
rect 4090 1038 4094 1041
rect 3990 952 3993 958
rect 3998 942 4001 948
rect 4006 932 4009 968
rect 4022 962 4025 978
rect 4062 972 4065 1018
rect 4070 992 4073 998
rect 4094 992 4097 1028
rect 4134 972 4137 1038
rect 4142 992 4145 1038
rect 4206 1031 4209 1058
rect 4238 1052 4241 1058
rect 4266 1048 4270 1051
rect 4218 1038 4225 1041
rect 4206 1028 4217 1031
rect 4098 968 4102 971
rect 3976 903 3978 907
rect 3982 903 3985 907
rect 3989 903 3992 907
rect 3710 742 3713 768
rect 3742 762 3745 768
rect 3750 752 3753 828
rect 3766 792 3769 848
rect 3862 792 3865 828
rect 3886 792 3889 818
rect 3894 802 3897 868
rect 3902 862 3905 868
rect 3934 862 3937 868
rect 3822 772 3825 778
rect 3854 772 3857 778
rect 3842 768 3846 771
rect 3874 768 3878 771
rect 3910 762 3913 858
rect 3930 848 3934 851
rect 3918 842 3921 848
rect 3942 842 3945 878
rect 3998 862 4001 918
rect 3974 852 3977 858
rect 3998 852 4001 858
rect 4006 852 4009 888
rect 4022 882 4025 928
rect 4014 862 4017 868
rect 3926 792 3929 798
rect 3934 772 3937 818
rect 3942 782 3945 838
rect 3958 792 3961 848
rect 4014 842 4017 848
rect 4022 842 4025 878
rect 4030 872 4033 948
rect 4038 932 4041 968
rect 4090 958 4094 961
rect 4066 948 4070 951
rect 4046 942 4049 948
rect 4054 892 4057 938
rect 4034 858 4046 861
rect 4062 852 4065 898
rect 4070 852 4073 908
rect 4078 902 4081 958
rect 4118 952 4121 958
rect 4094 942 4097 948
rect 4126 942 4129 948
rect 4078 862 4081 868
rect 4042 838 4046 841
rect 3966 832 3969 838
rect 4006 792 4009 838
rect 4038 792 4041 828
rect 4062 811 4065 848
rect 4086 842 4089 928
rect 4118 882 4121 888
rect 4094 872 4097 878
rect 4118 862 4121 868
rect 4126 852 4129 898
rect 4150 892 4153 1028
rect 4206 992 4209 1018
rect 4214 1001 4217 1028
rect 4222 1022 4225 1038
rect 4230 1032 4233 1048
rect 4242 1038 4246 1041
rect 4214 998 4225 1001
rect 4222 992 4225 998
rect 4246 972 4249 1038
rect 4270 992 4273 1028
rect 4286 992 4289 1058
rect 4234 968 4238 971
rect 4170 948 4174 951
rect 4182 922 4185 958
rect 4158 902 4161 918
rect 4182 892 4185 908
rect 4190 892 4193 948
rect 4198 932 4201 968
rect 4210 958 4214 961
rect 4250 958 4254 961
rect 4226 948 4230 951
rect 4222 942 4225 948
rect 4198 892 4201 918
rect 4222 892 4225 928
rect 4162 878 4166 881
rect 4134 862 4137 868
rect 4142 852 4145 868
rect 4110 832 4113 838
rect 4062 808 4073 811
rect 4062 792 4065 798
rect 3922 768 3926 771
rect 3954 768 3958 771
rect 3794 758 3798 761
rect 3834 758 3838 761
rect 3930 758 3934 761
rect 3806 752 3809 758
rect 3818 748 3822 751
rect 3850 748 3854 751
rect 3914 748 3918 751
rect 3946 748 3950 751
rect 3678 682 3681 718
rect 3678 672 3681 678
rect 3686 672 3689 678
rect 3694 672 3697 698
rect 3686 661 3689 668
rect 3678 658 3689 661
rect 3614 562 3617 648
rect 3646 642 3649 648
rect 3614 542 3617 558
rect 3614 482 3617 528
rect 3630 472 3633 638
rect 3638 592 3641 608
rect 3654 582 3657 648
rect 3678 612 3681 658
rect 3650 548 3654 551
rect 3642 538 3646 541
rect 3646 532 3649 538
rect 3630 462 3633 468
rect 3638 462 3641 498
rect 3646 472 3649 488
rect 3670 462 3673 518
rect 3594 448 3598 451
rect 3646 442 3649 458
rect 3678 452 3681 578
rect 3686 542 3689 618
rect 3702 572 3705 718
rect 3718 682 3721 738
rect 3718 672 3721 678
rect 3726 662 3729 748
rect 3786 738 3790 741
rect 3742 732 3745 738
rect 3798 732 3801 738
rect 3766 702 3769 718
rect 3742 692 3745 698
rect 3782 682 3785 728
rect 3750 672 3753 678
rect 3774 672 3777 678
rect 3798 672 3801 698
rect 3846 672 3849 698
rect 3854 682 3857 738
rect 3886 732 3889 748
rect 3910 692 3913 728
rect 3834 668 3838 671
rect 3806 662 3809 668
rect 3722 658 3726 661
rect 3754 658 3758 661
rect 3774 652 3777 658
rect 3746 648 3750 651
rect 3710 612 3713 618
rect 3714 588 3718 591
rect 3790 562 3793 618
rect 3722 558 3726 561
rect 3778 558 3782 561
rect 3746 548 3750 551
rect 3798 542 3801 658
rect 3822 652 3825 658
rect 3846 652 3849 658
rect 3830 642 3833 648
rect 3806 622 3809 628
rect 3806 562 3809 568
rect 3830 562 3833 638
rect 3746 538 3750 541
rect 3646 382 3649 438
rect 3654 402 3657 418
rect 3630 362 3633 378
rect 3638 352 3641 358
rect 3662 352 3665 448
rect 3678 392 3681 448
rect 3686 382 3689 538
rect 3822 532 3825 538
rect 3846 532 3849 538
rect 3702 472 3705 478
rect 3694 462 3697 468
rect 3670 362 3673 378
rect 3610 348 3614 351
rect 3674 338 3678 341
rect 3606 322 3609 338
rect 3646 322 3649 328
rect 3502 292 3505 298
rect 3526 282 3529 288
rect 3494 272 3497 278
rect 3518 262 3521 278
rect 3558 272 3561 298
rect 3574 272 3577 278
rect 3562 268 3566 271
rect 3542 262 3545 268
rect 3554 258 3558 261
rect 3566 252 3569 258
rect 3582 252 3585 288
rect 3590 262 3593 308
rect 3634 288 3638 291
rect 3606 282 3609 288
rect 3646 282 3649 318
rect 3618 278 3622 281
rect 3598 272 3601 278
rect 3598 252 3601 268
rect 3614 262 3617 278
rect 3662 272 3665 288
rect 3678 272 3681 318
rect 3694 282 3697 458
rect 3710 392 3713 468
rect 3726 422 3729 458
rect 3718 362 3721 418
rect 3718 351 3721 358
rect 3714 348 3721 351
rect 3734 342 3737 518
rect 3766 482 3769 518
rect 3790 492 3793 518
rect 3814 512 3817 518
rect 3746 468 3750 471
rect 3762 468 3766 471
rect 3786 468 3790 471
rect 3798 462 3801 508
rect 3814 471 3817 508
rect 3814 468 3822 471
rect 3778 458 3782 461
rect 3818 458 3822 461
rect 3818 448 3822 451
rect 3774 352 3777 418
rect 3798 412 3801 418
rect 3810 368 3814 371
rect 3830 361 3833 518
rect 3854 482 3857 678
rect 3862 662 3865 678
rect 3870 672 3873 678
rect 3878 662 3881 668
rect 3886 662 3889 678
rect 3898 648 3902 651
rect 3894 562 3897 618
rect 3910 572 3913 658
rect 3918 572 3921 638
rect 3926 592 3929 748
rect 3934 592 3937 648
rect 3942 572 3945 658
rect 3958 641 3961 768
rect 3966 712 3969 758
rect 3990 752 3993 788
rect 4002 768 4006 771
rect 3976 703 3978 707
rect 3982 703 3985 707
rect 3989 703 3992 707
rect 3998 692 4001 758
rect 4014 722 4017 758
rect 4022 752 4025 788
rect 4050 768 4054 771
rect 4030 732 4033 768
rect 4070 762 4073 808
rect 4134 792 4137 838
rect 4158 822 4161 868
rect 4166 852 4169 858
rect 4062 742 4065 748
rect 3998 642 4001 658
rect 4006 652 4009 658
rect 4014 652 4017 688
rect 4022 662 4025 668
rect 4042 658 4046 661
rect 4058 658 4062 661
rect 4070 652 4073 758
rect 4102 752 4105 768
rect 4110 752 4113 758
rect 4118 752 4121 758
rect 4126 732 4129 768
rect 4166 742 4169 748
rect 4086 672 4089 718
rect 4078 642 4081 648
rect 4086 642 4089 658
rect 4094 642 4097 728
rect 4150 681 4153 718
rect 4158 692 4161 708
rect 4174 682 4177 878
rect 4190 872 4193 878
rect 4206 862 4209 868
rect 4234 858 4238 861
rect 4190 792 4193 818
rect 4230 792 4233 818
rect 4238 782 4241 848
rect 4226 768 4230 771
rect 4150 678 4161 681
rect 4170 678 4174 681
rect 4126 672 4129 678
rect 4146 668 4150 671
rect 4102 662 4105 668
rect 4122 658 4126 661
rect 3954 638 3961 641
rect 3986 638 3990 641
rect 3966 592 3969 638
rect 3974 632 3977 638
rect 4006 592 4009 638
rect 4022 592 4025 638
rect 4030 582 4033 638
rect 4054 632 4057 638
rect 4062 632 4065 638
rect 4070 592 4073 638
rect 4030 572 4033 578
rect 3874 558 3878 561
rect 3902 552 3905 558
rect 3910 552 3913 568
rect 3918 562 3921 568
rect 3926 558 3934 561
rect 3882 538 3886 541
rect 3842 478 3846 481
rect 3862 472 3865 518
rect 3874 478 3878 481
rect 3894 472 3897 518
rect 3914 478 3918 481
rect 3882 468 3886 471
rect 3838 452 3841 458
rect 3854 402 3857 458
rect 3854 372 3857 378
rect 3862 372 3865 468
rect 3822 358 3833 361
rect 3838 362 3841 368
rect 3870 362 3873 458
rect 3722 338 3726 341
rect 3746 338 3750 341
rect 3730 328 3734 331
rect 3406 152 3409 178
rect 3414 142 3417 148
rect 3426 138 3430 141
rect 3434 128 3438 131
rect 3282 88 3289 91
rect 3346 88 3350 91
rect 3254 72 3257 78
rect 3162 68 3166 71
rect 3210 68 3214 71
rect 3198 62 3201 68
rect 3334 62 3337 68
rect 2778 58 2782 61
rect 2938 58 2942 61
rect 3170 58 3174 61
rect 3186 58 3190 61
rect 3242 58 3246 61
rect 2742 52 2745 58
rect 2294 -18 2297 28
rect 2310 22 2313 48
rect 2310 -18 2313 18
rect 2398 12 2401 48
rect 2574 22 2577 50
rect 2642 48 2646 51
rect 2666 48 2670 51
rect 2934 22 2937 48
rect 3126 31 3129 50
rect 3190 42 3193 48
rect 3230 32 3233 58
rect 3266 48 3270 51
rect 3374 32 3377 118
rect 3430 82 3433 108
rect 3454 102 3457 218
rect 3472 203 3474 207
rect 3478 203 3481 207
rect 3485 203 3488 207
rect 3466 168 3470 171
rect 3502 152 3505 248
rect 3446 72 3449 78
rect 3502 62 3505 148
rect 3542 132 3545 218
rect 3558 142 3561 208
rect 3606 162 3609 188
rect 3622 172 3625 268
rect 3678 262 3681 268
rect 3702 262 3705 318
rect 3734 302 3737 328
rect 3718 262 3721 278
rect 3758 272 3761 318
rect 3766 292 3769 328
rect 3774 322 3777 348
rect 3822 342 3825 358
rect 3834 348 3838 351
rect 3846 331 3849 358
rect 3878 351 3881 368
rect 3886 361 3889 468
rect 3894 462 3897 468
rect 3886 358 3897 361
rect 3878 348 3886 351
rect 3854 342 3857 348
rect 3894 342 3897 358
rect 3902 352 3905 458
rect 3926 432 3929 558
rect 3942 552 3945 568
rect 3950 562 3953 568
rect 3934 462 3937 468
rect 3942 462 3945 478
rect 3958 462 3961 568
rect 3966 562 3969 568
rect 3942 381 3945 458
rect 3950 442 3953 448
rect 3966 442 3969 558
rect 3982 552 3985 558
rect 3990 552 3993 568
rect 3976 503 3978 507
rect 3982 503 3985 507
rect 3989 503 3992 507
rect 3998 492 4001 508
rect 4014 492 4017 558
rect 4026 548 4030 551
rect 4002 468 4006 471
rect 3986 448 3990 451
rect 3966 432 3969 438
rect 3934 378 3945 381
rect 3934 352 3937 378
rect 3942 352 3945 368
rect 3982 352 3985 418
rect 4006 392 4009 468
rect 4022 462 4025 548
rect 4038 481 4041 578
rect 4062 572 4065 578
rect 4086 572 4089 638
rect 4118 592 4121 638
rect 4134 622 4137 648
rect 4142 632 4145 658
rect 4102 582 4105 588
rect 4094 572 4097 578
rect 4158 572 4161 678
rect 4166 642 4169 668
rect 4098 568 4102 571
rect 4130 568 4134 571
rect 4174 562 4177 648
rect 4182 592 4185 768
rect 4198 752 4201 758
rect 4190 722 4193 748
rect 4206 692 4209 758
rect 4218 748 4222 751
rect 4214 692 4217 718
rect 4198 662 4201 668
rect 4218 658 4222 661
rect 4206 622 4209 648
rect 4214 592 4217 638
rect 4230 572 4233 768
rect 4238 752 4241 778
rect 4246 692 4249 938
rect 4254 902 4257 948
rect 4274 938 4278 941
rect 4254 882 4257 888
rect 4270 862 4273 928
rect 4286 922 4289 948
rect 4294 911 4297 1068
rect 4310 1061 4313 1068
rect 4326 1062 4329 1128
rect 4358 1102 4361 1148
rect 4342 1092 4345 1098
rect 4374 1092 4377 1168
rect 4310 1058 4318 1061
rect 4302 962 4305 1048
rect 4310 952 4313 1058
rect 4326 932 4329 1058
rect 4286 908 4297 911
rect 4278 892 4281 908
rect 4270 852 4273 858
rect 4286 851 4289 908
rect 4318 882 4321 898
rect 4318 862 4321 878
rect 4282 848 4289 851
rect 4294 842 4297 858
rect 4302 852 4305 858
rect 4310 852 4313 858
rect 4326 852 4329 918
rect 4342 892 4345 1068
rect 4358 1062 4361 1088
rect 4358 942 4361 1058
rect 4374 952 4377 1078
rect 4350 882 4353 918
rect 4346 838 4350 841
rect 4286 822 4289 838
rect 4326 832 4329 838
rect 4334 832 4337 838
rect 4358 822 4361 858
rect 4366 842 4369 848
rect 4278 772 4281 778
rect 4302 762 4305 808
rect 4326 792 4329 818
rect 4314 768 4318 771
rect 4374 762 4377 948
rect 4306 748 4310 751
rect 4254 742 4257 748
rect 4294 742 4297 748
rect 4226 568 4230 571
rect 4190 562 4193 568
rect 4074 558 4078 561
rect 4106 558 4110 561
rect 4138 558 4142 561
rect 4178 558 4182 561
rect 4046 522 4049 558
rect 4166 552 4169 558
rect 4058 548 4062 551
rect 4082 548 4086 551
rect 4114 548 4118 551
rect 4146 548 4150 551
rect 4178 548 4182 551
rect 4030 478 4041 481
rect 4014 362 4017 448
rect 4030 442 4033 478
rect 4038 462 4041 468
rect 3866 338 3870 341
rect 3906 338 3910 341
rect 3846 328 3857 331
rect 3790 322 3793 328
rect 3806 292 3809 328
rect 3794 288 3798 291
rect 3806 282 3809 288
rect 3794 268 3801 271
rect 3726 262 3729 268
rect 3754 258 3758 261
rect 3634 248 3638 251
rect 3638 192 3641 218
rect 3654 192 3657 218
rect 3634 188 3638 191
rect 3614 152 3617 158
rect 3534 72 3537 88
rect 3550 62 3553 68
rect 3558 62 3561 118
rect 3606 92 3609 98
rect 3574 52 3577 88
rect 3582 62 3585 88
rect 3606 82 3609 88
rect 3614 72 3617 138
rect 3662 122 3665 258
rect 3714 248 3718 251
rect 3702 222 3705 248
rect 3726 232 3729 258
rect 3738 248 3742 251
rect 3766 232 3769 268
rect 3798 262 3801 268
rect 3814 270 3817 298
rect 3854 272 3857 328
rect 3870 281 3873 318
rect 3862 278 3873 281
rect 3750 212 3753 218
rect 3634 78 3638 81
rect 3614 62 3617 68
rect 3638 52 3641 68
rect 3646 62 3649 78
rect 3670 62 3673 158
rect 3678 72 3681 198
rect 3718 132 3721 208
rect 3774 192 3777 258
rect 3766 160 3769 179
rect 3734 152 3737 158
rect 3734 132 3737 138
rect 3702 92 3705 98
rect 3718 91 3721 118
rect 3774 101 3777 148
rect 3790 122 3793 248
rect 3806 142 3809 268
rect 3814 182 3817 266
rect 3862 262 3865 278
rect 3886 272 3889 318
rect 3894 272 3897 338
rect 3926 332 3929 338
rect 3918 302 3921 318
rect 3934 282 3937 328
rect 3922 278 3929 281
rect 3926 272 3929 278
rect 3934 272 3937 278
rect 3950 272 3953 338
rect 3966 332 3969 338
rect 3958 311 3961 318
rect 3958 308 3966 311
rect 3976 303 3978 307
rect 3982 303 3985 307
rect 3989 303 3992 307
rect 3982 282 3985 288
rect 3998 272 4001 338
rect 4046 292 4049 498
rect 4062 472 4065 478
rect 4102 462 4105 468
rect 4126 462 4129 548
rect 4190 492 4193 548
rect 4206 532 4209 558
rect 4214 532 4217 548
rect 4206 482 4209 518
rect 4202 478 4206 481
rect 4158 472 4161 478
rect 4182 472 4185 478
rect 4174 462 4177 468
rect 4214 462 4217 528
rect 4238 522 4241 678
rect 4334 672 4337 758
rect 4390 752 4393 1178
rect 4362 748 4366 751
rect 4342 722 4345 728
rect 4270 668 4278 671
rect 4254 592 4257 668
rect 4270 661 4273 668
rect 4334 662 4337 668
rect 4266 658 4273 661
rect 4314 658 4318 661
rect 4266 648 4270 651
rect 4246 572 4249 578
rect 4262 562 4265 618
rect 4270 612 4273 648
rect 4270 562 4273 598
rect 4278 592 4281 658
rect 4298 648 4302 651
rect 4342 642 4345 718
rect 4374 672 4377 718
rect 4386 678 4390 681
rect 4350 662 4353 668
rect 4290 638 4294 641
rect 4322 638 4326 641
rect 4310 632 4313 638
rect 4358 592 4361 668
rect 4370 658 4377 661
rect 4282 568 4286 571
rect 4314 568 4318 571
rect 4366 562 4369 608
rect 4374 592 4377 658
rect 4378 568 4382 571
rect 4258 558 4262 561
rect 4330 558 4334 561
rect 4270 548 4278 551
rect 4242 488 4246 491
rect 4222 462 4225 468
rect 4246 462 4249 468
rect 4254 462 4257 548
rect 4286 538 4294 541
rect 4286 492 4289 538
rect 4302 512 4305 558
rect 4314 548 4318 551
rect 4270 462 4273 488
rect 4282 468 4286 471
rect 4058 458 4062 461
rect 4090 458 4094 461
rect 4154 458 4158 461
rect 4082 448 4086 451
rect 4130 448 4134 451
rect 4170 448 4174 451
rect 4054 442 4057 448
rect 4070 402 4073 448
rect 4114 438 4118 441
rect 4146 438 4150 441
rect 4094 432 4097 438
rect 4126 432 4129 438
rect 4182 392 4185 458
rect 4206 422 4209 448
rect 4226 438 4230 441
rect 4214 392 4217 428
rect 4246 392 4249 438
rect 4262 402 4265 448
rect 4278 392 4281 458
rect 4294 432 4297 478
rect 4310 472 4313 478
rect 4326 452 4329 558
rect 4346 548 4350 551
rect 4342 462 4345 528
rect 4306 448 4310 451
rect 4338 448 4342 451
rect 4330 438 4334 441
rect 4310 392 4313 438
rect 4318 432 4321 438
rect 4342 422 4345 428
rect 4358 392 4361 548
rect 4374 492 4377 548
rect 4370 458 4374 461
rect 4150 362 4153 388
rect 4194 368 4198 371
rect 4226 368 4230 371
rect 4258 368 4262 371
rect 4270 362 4273 378
rect 4290 368 4294 371
rect 4322 368 4326 371
rect 4354 368 4358 371
rect 4170 358 4174 361
rect 4202 358 4206 361
rect 4234 358 4238 361
rect 4298 358 4302 361
rect 4278 352 4281 358
rect 4186 348 4190 351
rect 4218 348 4222 351
rect 4250 348 4254 351
rect 4306 348 4310 351
rect 4102 342 4105 348
rect 4086 332 4089 338
rect 4102 272 4105 278
rect 4010 268 4014 271
rect 4082 268 4086 271
rect 3870 262 3873 268
rect 3998 262 4001 268
rect 3890 258 3894 261
rect 3906 258 3910 261
rect 3938 258 3942 261
rect 4018 258 4022 261
rect 4042 258 4046 261
rect 3830 232 3833 248
rect 3846 242 3849 258
rect 3902 232 3905 248
rect 3918 242 3921 258
rect 3954 248 3958 251
rect 4006 251 4009 258
rect 3998 248 4009 251
rect 3870 222 3873 228
rect 3894 182 3897 198
rect 3834 158 3838 161
rect 3814 152 3817 158
rect 3854 152 3857 158
rect 3838 142 3841 148
rect 3846 142 3849 148
rect 3862 132 3865 178
rect 3878 152 3881 158
rect 3894 152 3897 178
rect 3922 158 3926 161
rect 3902 152 3905 158
rect 3934 152 3937 158
rect 3918 142 3921 148
rect 3926 142 3929 148
rect 3958 142 3961 248
rect 3978 238 3982 241
rect 3998 232 4001 248
rect 4038 242 4041 248
rect 3998 192 4001 228
rect 4030 192 4033 218
rect 4046 212 4049 248
rect 3966 152 3969 178
rect 4062 172 4065 258
rect 4070 232 4073 268
rect 4134 262 4137 348
rect 4334 312 4337 358
rect 4346 348 4350 351
rect 4350 292 4353 328
rect 4366 322 4369 448
rect 4378 438 4382 441
rect 4274 288 4278 291
rect 4198 282 4201 288
rect 4182 272 4185 278
rect 4078 252 4081 258
rect 4110 232 4113 258
rect 4086 202 4089 218
rect 3970 148 3974 151
rect 4010 148 4014 151
rect 3882 138 3886 141
rect 3942 132 3945 138
rect 3950 132 3953 138
rect 3834 118 3838 121
rect 3714 88 3721 91
rect 3766 98 3777 101
rect 3710 82 3713 88
rect 3722 68 3725 71
rect 3686 62 3689 68
rect 3694 52 3697 68
rect 3766 62 3769 98
rect 3806 82 3809 98
rect 3902 92 3905 98
rect 3966 92 3969 138
rect 3976 103 3978 107
rect 3982 103 3985 107
rect 3989 103 3992 107
rect 4038 92 4041 158
rect 4038 82 4041 88
rect 3822 72 3825 78
rect 3958 72 3961 78
rect 3878 62 3881 68
rect 3966 62 3969 68
rect 4054 62 4057 108
rect 4070 72 4073 148
rect 4110 132 4113 168
rect 4126 152 4129 258
rect 4150 231 4153 250
rect 4174 162 4177 188
rect 4206 172 4209 178
rect 4126 132 4129 138
rect 4086 92 4089 108
rect 4102 62 4105 68
rect 4118 62 4121 68
rect 4134 62 4137 108
rect 4174 92 4177 108
rect 4170 78 4174 81
rect 4142 72 4145 78
rect 4150 62 4153 78
rect 4166 72 4169 78
rect 4190 62 4193 138
rect 4214 92 4217 208
rect 4262 162 4265 278
rect 4286 272 4289 278
rect 4286 192 4289 258
rect 4270 162 4273 178
rect 4262 142 4265 158
rect 4286 152 4289 168
rect 4262 92 4265 118
rect 4294 92 4297 228
rect 4334 192 4337 258
rect 4366 192 4369 308
rect 4318 152 4321 158
rect 4302 142 4305 148
rect 4302 122 4305 128
rect 4310 122 4313 128
rect 4198 72 4201 88
rect 4206 62 4209 68
rect 4246 62 4249 78
rect 4278 62 4281 68
rect 3610 48 3614 51
rect 4310 52 4313 118
rect 4318 62 4321 68
rect 3494 22 3497 48
rect 3654 42 3657 48
rect 3670 42 3673 48
rect 3854 22 3857 50
rect 4162 48 4166 51
rect 4174 42 4177 48
rect 4326 42 4329 158
rect 4334 92 4337 178
rect 4390 172 4393 618
rect 4362 158 4366 161
rect 4350 112 4353 148
rect 4374 132 4377 138
rect 4358 92 4361 98
rect 4338 58 4342 61
rect 4070 12 4073 18
rect 2398 -18 2401 8
rect 2440 3 2442 7
rect 2446 3 2449 7
rect 2453 3 2456 7
rect 2566 -18 2569 8
rect 2638 -18 2641 8
rect 2750 -18 2753 8
rect 3472 3 3474 7
rect 3478 3 3481 7
rect 3485 3 3488 7
rect 4054 -18 4057 8
rect 1358 -19 1362 -18
rect 1350 -22 1362 -19
rect 1374 -22 1378 -18
rect 1438 -22 1442 -18
rect 1598 -22 1602 -18
rect 2022 -22 2026 -18
rect 2134 -22 2138 -18
rect 2150 -22 2154 -18
rect 2166 -22 2170 -18
rect 2270 -22 2274 -18
rect 2294 -22 2298 -18
rect 2310 -22 2314 -18
rect 2398 -22 2402 -18
rect 2566 -22 2570 -18
rect 2638 -22 2642 -18
rect 2750 -22 2754 -18
rect 3694 -22 3698 -18
rect 4054 -22 4058 -18
<< m3contact >>
rect 898 3103 902 3107
rect 905 3103 909 3107
rect 1134 3098 1138 3102
rect 1158 3098 1162 3102
rect 1198 3098 1202 3102
rect 1254 3098 1258 3102
rect 1270 3098 1274 3102
rect 1358 3098 1362 3102
rect 1470 3098 1474 3102
rect 654 3088 658 3092
rect 678 3088 682 3092
rect 686 3088 690 3092
rect 838 3088 842 3092
rect 214 3078 218 3082
rect 438 3078 442 3082
rect 566 3078 570 3082
rect 598 3078 602 3082
rect 622 3078 626 3082
rect 230 3068 234 3072
rect 454 3068 458 3072
rect 558 3068 562 3072
rect 614 3068 618 3072
rect 30 3058 34 3062
rect 78 3058 82 3062
rect 230 3058 234 3062
rect 318 3058 322 3062
rect 566 3058 570 3062
rect 582 3058 586 3062
rect 622 3058 626 3062
rect 6 3018 10 3022
rect 14 2778 18 2782
rect 134 2998 138 3002
rect 214 3048 218 3052
rect 182 3038 186 3042
rect 310 3048 314 3052
rect 262 2998 266 3002
rect 174 2938 178 2942
rect 62 2908 66 2912
rect 110 2908 114 2912
rect 102 2878 106 2882
rect 94 2838 98 2842
rect 158 2828 162 2832
rect 22 2768 26 2772
rect 70 2778 74 2782
rect 38 2758 42 2762
rect 262 2898 266 2902
rect 278 2878 282 2882
rect 238 2858 242 2862
rect 214 2828 218 2832
rect 246 2828 250 2832
rect 262 2858 266 2862
rect 334 3038 338 3042
rect 382 3048 386 3052
rect 542 3028 546 3032
rect 394 3003 398 3007
rect 401 3003 405 3007
rect 350 2988 354 2992
rect 478 2988 482 2992
rect 350 2948 354 2952
rect 374 2948 378 2952
rect 382 2948 386 2952
rect 430 2948 434 2952
rect 350 2938 354 2942
rect 542 2938 546 2942
rect 422 2928 426 2932
rect 438 2928 442 2932
rect 414 2918 418 2922
rect 358 2898 362 2902
rect 342 2878 346 2882
rect 302 2828 306 2832
rect 254 2808 258 2812
rect 198 2788 202 2792
rect 174 2778 178 2782
rect 86 2768 90 2772
rect 326 2788 330 2792
rect 102 2758 106 2762
rect 158 2758 162 2762
rect 30 2748 34 2752
rect 166 2748 170 2752
rect 38 2738 42 2742
rect 54 2738 58 2742
rect 86 2738 90 2742
rect 142 2738 146 2742
rect 78 2728 82 2732
rect 102 2728 106 2732
rect 182 2728 186 2732
rect 118 2718 122 2722
rect 174 2718 178 2722
rect 94 2708 98 2712
rect 62 2698 66 2702
rect 70 2678 74 2682
rect 270 2748 274 2752
rect 246 2738 250 2742
rect 222 2718 226 2722
rect 198 2708 202 2712
rect 206 2708 210 2712
rect 198 2688 202 2692
rect 142 2668 146 2672
rect 190 2668 194 2672
rect 86 2618 90 2622
rect 38 2598 42 2602
rect 94 2588 98 2592
rect 30 2568 34 2572
rect 6 2548 10 2552
rect 118 2558 122 2562
rect 118 2548 122 2552
rect 174 2648 178 2652
rect 230 2688 234 2692
rect 222 2678 226 2682
rect 286 2738 290 2742
rect 278 2728 282 2732
rect 310 2748 314 2752
rect 318 2738 322 2742
rect 350 2808 354 2812
rect 342 2768 346 2772
rect 326 2718 330 2722
rect 302 2708 306 2712
rect 262 2678 266 2682
rect 318 2678 322 2682
rect 238 2668 242 2672
rect 394 2803 398 2807
rect 401 2803 405 2807
rect 574 2928 578 2932
rect 558 2918 562 2922
rect 430 2888 434 2892
rect 478 2868 482 2872
rect 518 2898 522 2902
rect 542 2898 546 2902
rect 566 2898 570 2902
rect 574 2878 578 2882
rect 550 2868 554 2872
rect 718 3078 722 3082
rect 798 3078 802 3082
rect 654 3068 658 3072
rect 790 3068 794 3072
rect 694 3058 698 3062
rect 630 3028 634 3032
rect 590 2978 594 2982
rect 622 2978 626 2982
rect 606 2948 610 2952
rect 614 2948 618 2952
rect 686 2968 690 2972
rect 654 2948 658 2952
rect 678 2948 682 2952
rect 670 2938 674 2942
rect 622 2928 626 2932
rect 646 2928 650 2932
rect 654 2918 658 2922
rect 662 2918 666 2922
rect 646 2908 650 2912
rect 646 2888 650 2892
rect 598 2878 602 2882
rect 590 2868 594 2872
rect 622 2868 626 2872
rect 502 2858 506 2862
rect 470 2818 474 2822
rect 438 2808 442 2812
rect 422 2788 426 2792
rect 462 2788 466 2792
rect 358 2778 362 2782
rect 462 2758 466 2762
rect 430 2728 434 2732
rect 414 2718 418 2722
rect 414 2708 418 2712
rect 382 2678 386 2682
rect 294 2668 298 2672
rect 334 2668 338 2672
rect 350 2668 354 2672
rect 214 2658 218 2662
rect 254 2658 258 2662
rect 278 2658 282 2662
rect 254 2648 258 2652
rect 214 2628 218 2632
rect 238 2628 242 2632
rect 262 2588 266 2592
rect 270 2588 274 2592
rect 214 2568 218 2572
rect 198 2558 202 2562
rect 230 2558 234 2562
rect 206 2548 210 2552
rect 246 2548 250 2552
rect 86 2538 90 2542
rect 150 2538 154 2542
rect 174 2538 178 2542
rect 190 2538 194 2542
rect 214 2538 218 2542
rect 270 2538 274 2542
rect 22 2528 26 2532
rect 230 2508 234 2512
rect 70 2498 74 2502
rect 110 2498 114 2502
rect 126 2498 130 2502
rect 166 2498 170 2502
rect 174 2498 178 2502
rect 214 2498 218 2502
rect 86 2488 90 2492
rect 190 2478 194 2482
rect 422 2698 426 2702
rect 438 2678 442 2682
rect 358 2658 362 2662
rect 374 2658 378 2662
rect 302 2648 306 2652
rect 414 2638 418 2642
rect 422 2608 426 2612
rect 394 2603 398 2607
rect 401 2603 405 2607
rect 358 2498 362 2502
rect 294 2488 298 2492
rect 390 2508 394 2512
rect 382 2488 386 2492
rect 310 2478 314 2482
rect 374 2478 378 2482
rect 238 2468 242 2472
rect 294 2458 298 2462
rect 414 2458 418 2462
rect 30 2450 34 2454
rect 366 2448 370 2452
rect 430 2528 434 2532
rect 478 2758 482 2762
rect 478 2688 482 2692
rect 486 2608 490 2612
rect 486 2598 490 2602
rect 470 2558 474 2562
rect 454 2508 458 2512
rect 502 2798 506 2802
rect 534 2798 538 2802
rect 526 2788 530 2792
rect 558 2858 562 2862
rect 582 2858 586 2862
rect 574 2838 578 2842
rect 550 2778 554 2782
rect 526 2758 530 2762
rect 534 2758 538 2762
rect 502 2748 506 2752
rect 510 2738 514 2742
rect 534 2738 538 2742
rect 518 2728 522 2732
rect 534 2728 538 2732
rect 630 2838 634 2842
rect 606 2818 610 2822
rect 574 2748 578 2752
rect 582 2748 586 2752
rect 574 2728 578 2732
rect 566 2718 570 2722
rect 558 2708 562 2712
rect 550 2698 554 2702
rect 566 2698 570 2702
rect 502 2658 506 2662
rect 526 2658 530 2662
rect 550 2658 554 2662
rect 526 2638 530 2642
rect 534 2638 538 2642
rect 542 2608 546 2612
rect 630 2758 634 2762
rect 606 2728 610 2732
rect 598 2668 602 2672
rect 574 2658 578 2662
rect 558 2648 562 2652
rect 566 2638 570 2642
rect 550 2598 554 2602
rect 510 2578 514 2582
rect 510 2568 514 2572
rect 526 2568 530 2572
rect 478 2538 482 2542
rect 486 2538 490 2542
rect 518 2538 522 2542
rect 542 2538 546 2542
rect 494 2528 498 2532
rect 590 2648 594 2652
rect 670 2898 674 2902
rect 662 2868 666 2872
rect 734 3058 738 3062
rect 1054 3078 1058 3082
rect 878 3068 882 3072
rect 950 3068 954 3072
rect 814 3058 818 3062
rect 838 3058 842 3062
rect 710 3048 714 3052
rect 830 3048 834 3052
rect 854 3048 858 3052
rect 726 3038 730 3042
rect 750 3038 754 3042
rect 702 3028 706 3032
rect 822 2978 826 2982
rect 878 2968 882 2972
rect 870 2958 874 2962
rect 766 2938 770 2942
rect 814 2938 818 2942
rect 830 2938 834 2942
rect 782 2928 786 2932
rect 742 2818 746 2822
rect 694 2798 698 2802
rect 686 2768 690 2772
rect 670 2758 674 2762
rect 718 2758 722 2762
rect 766 2858 770 2862
rect 854 2908 858 2912
rect 838 2898 842 2902
rect 958 3048 962 3052
rect 942 3038 946 3042
rect 982 3038 986 3042
rect 926 3028 930 3032
rect 974 2968 978 2972
rect 902 2918 906 2922
rect 942 2928 946 2932
rect 950 2928 954 2932
rect 958 2918 962 2922
rect 926 2908 930 2912
rect 950 2908 954 2912
rect 974 2908 978 2912
rect 898 2903 902 2907
rect 905 2903 909 2907
rect 926 2898 930 2902
rect 942 2888 946 2892
rect 918 2878 922 2882
rect 806 2798 810 2802
rect 758 2758 762 2762
rect 638 2748 642 2752
rect 734 2748 738 2752
rect 750 2748 754 2752
rect 798 2748 802 2752
rect 742 2738 746 2742
rect 694 2728 698 2732
rect 718 2728 722 2732
rect 622 2648 626 2652
rect 614 2628 618 2632
rect 646 2648 650 2652
rect 638 2608 642 2612
rect 782 2728 786 2732
rect 806 2728 810 2732
rect 774 2718 778 2722
rect 806 2718 810 2722
rect 750 2708 754 2712
rect 678 2698 682 2702
rect 670 2658 674 2662
rect 662 2618 666 2622
rect 598 2578 602 2582
rect 590 2568 594 2572
rect 630 2568 634 2572
rect 598 2548 602 2552
rect 590 2538 594 2542
rect 566 2528 570 2532
rect 582 2528 586 2532
rect 486 2508 490 2512
rect 542 2508 546 2512
rect 550 2508 554 2512
rect 566 2508 570 2512
rect 502 2478 506 2482
rect 422 2448 426 2452
rect 414 2438 418 2442
rect 438 2418 442 2422
rect 394 2403 398 2407
rect 401 2403 405 2407
rect 358 2358 362 2362
rect 134 2348 138 2352
rect 190 2348 194 2352
rect 222 2348 226 2352
rect 286 2348 290 2352
rect 30 2338 34 2342
rect 214 2338 218 2342
rect 118 2318 122 2322
rect 22 2308 26 2312
rect 174 2288 178 2292
rect 190 2288 194 2292
rect 62 2278 66 2282
rect 30 2268 34 2272
rect 38 2268 42 2272
rect 478 2428 482 2432
rect 574 2488 578 2492
rect 606 2508 610 2512
rect 622 2488 626 2492
rect 550 2478 554 2482
rect 590 2478 594 2482
rect 542 2458 546 2462
rect 510 2448 514 2452
rect 526 2418 530 2422
rect 646 2528 650 2532
rect 638 2488 642 2492
rect 646 2478 650 2482
rect 630 2468 634 2472
rect 614 2458 618 2462
rect 614 2448 618 2452
rect 574 2418 578 2422
rect 622 2418 626 2422
rect 494 2408 498 2412
rect 558 2408 562 2412
rect 614 2348 618 2352
rect 430 2338 434 2342
rect 470 2338 474 2342
rect 566 2338 570 2342
rect 342 2328 346 2332
rect 262 2278 266 2282
rect 6 2258 10 2262
rect 22 2258 26 2262
rect 38 2248 42 2252
rect 54 2218 58 2222
rect 6 2178 10 2182
rect 54 2178 58 2182
rect 30 2158 34 2162
rect 70 2158 74 2162
rect 422 2258 426 2262
rect 366 2238 370 2242
rect 394 2203 398 2207
rect 401 2203 405 2207
rect 254 2188 258 2192
rect 270 2188 274 2192
rect 318 2188 322 2192
rect 310 2168 314 2172
rect 262 2158 266 2162
rect 30 2148 34 2152
rect 54 2148 58 2152
rect 78 2148 82 2152
rect 182 2148 186 2152
rect 302 2148 306 2152
rect 166 2138 170 2142
rect 46 2118 50 2122
rect 30 2068 34 2072
rect 182 2098 186 2102
rect 166 2088 170 2092
rect 62 2068 66 2072
rect 78 2068 82 2072
rect 342 2148 346 2152
rect 334 2128 338 2132
rect 294 2118 298 2122
rect 334 2088 338 2092
rect 286 2078 290 2082
rect 462 2258 466 2262
rect 414 2108 418 2112
rect 550 2308 554 2312
rect 534 2298 538 2302
rect 566 2298 570 2302
rect 654 2468 658 2472
rect 878 2858 882 2862
rect 894 2858 898 2862
rect 878 2848 882 2852
rect 822 2758 826 2762
rect 838 2758 842 2762
rect 870 2808 874 2812
rect 862 2768 866 2772
rect 870 2768 874 2772
rect 830 2748 834 2752
rect 854 2748 858 2752
rect 870 2748 874 2752
rect 862 2738 866 2742
rect 830 2728 834 2732
rect 854 2728 858 2732
rect 814 2698 818 2702
rect 854 2708 858 2712
rect 710 2678 714 2682
rect 814 2668 818 2672
rect 846 2688 850 2692
rect 854 2688 858 2692
rect 846 2678 850 2682
rect 870 2718 874 2722
rect 910 2758 914 2762
rect 1174 3058 1178 3062
rect 1286 3058 1290 3062
rect 1110 3048 1114 3052
rect 1134 3038 1138 3042
rect 1038 3028 1042 3032
rect 1174 3038 1178 3042
rect 1270 3038 1274 3042
rect 1030 2988 1034 2992
rect 1150 2988 1154 2992
rect 990 2958 994 2962
rect 1182 2988 1186 2992
rect 1174 2960 1178 2962
rect 1174 2958 1178 2960
rect 1006 2948 1010 2952
rect 998 2938 1002 2942
rect 1086 2938 1090 2942
rect 1046 2928 1050 2932
rect 1014 2888 1018 2892
rect 1078 2908 1082 2912
rect 1038 2878 1042 2882
rect 1062 2878 1066 2882
rect 966 2868 970 2872
rect 926 2838 930 2842
rect 966 2858 970 2862
rect 894 2748 898 2752
rect 918 2748 922 2752
rect 910 2728 914 2732
rect 886 2718 890 2722
rect 870 2688 874 2692
rect 726 2658 730 2662
rect 854 2648 858 2652
rect 790 2588 794 2592
rect 830 2558 834 2562
rect 726 2548 730 2552
rect 790 2498 794 2502
rect 830 2548 834 2552
rect 862 2548 866 2552
rect 898 2703 902 2707
rect 905 2703 909 2707
rect 894 2688 898 2692
rect 950 2768 954 2772
rect 982 2838 986 2842
rect 1054 2858 1058 2862
rect 1070 2858 1074 2862
rect 990 2768 994 2772
rect 1014 2768 1018 2772
rect 966 2738 970 2742
rect 974 2738 978 2742
rect 982 2728 986 2732
rect 998 2748 1002 2752
rect 1022 2748 1026 2752
rect 1046 2748 1050 2752
rect 1054 2748 1058 2752
rect 1006 2738 1010 2742
rect 950 2718 954 2722
rect 990 2718 994 2722
rect 1022 2718 1026 2722
rect 942 2678 946 2682
rect 918 2668 922 2672
rect 1046 2708 1050 2712
rect 1054 2678 1058 2682
rect 894 2648 898 2652
rect 878 2598 882 2602
rect 966 2568 970 2572
rect 950 2548 954 2552
rect 838 2538 842 2542
rect 870 2538 874 2542
rect 898 2503 902 2507
rect 905 2503 909 2507
rect 814 2488 818 2492
rect 926 2488 930 2492
rect 1142 2898 1146 2902
rect 1342 2978 1346 2982
rect 1238 2958 1242 2962
rect 1278 2928 1282 2932
rect 1294 2918 1298 2922
rect 1542 3068 1546 3072
rect 1534 3018 1538 3022
rect 1418 3003 1422 3007
rect 1425 3003 1429 3007
rect 1398 2988 1402 2992
rect 1406 2948 1410 2952
rect 1390 2928 1394 2932
rect 1270 2898 1274 2902
rect 1358 2898 1362 2902
rect 1206 2868 1210 2872
rect 1126 2838 1130 2842
rect 1254 2858 1258 2862
rect 1198 2828 1202 2832
rect 1182 2808 1186 2812
rect 1126 2798 1130 2802
rect 1150 2798 1154 2802
rect 1150 2788 1154 2792
rect 1166 2728 1170 2732
rect 1166 2718 1170 2722
rect 1142 2708 1146 2712
rect 1150 2698 1154 2702
rect 1182 2708 1186 2712
rect 1222 2808 1226 2812
rect 1246 2808 1250 2812
rect 1206 2748 1210 2752
rect 1214 2728 1218 2732
rect 1206 2718 1210 2722
rect 1214 2668 1218 2672
rect 1070 2608 1074 2612
rect 1046 2598 1050 2602
rect 1038 2498 1042 2502
rect 966 2478 970 2482
rect 990 2478 994 2482
rect 1006 2478 1010 2482
rect 742 2458 746 2462
rect 726 2438 730 2442
rect 726 2418 730 2422
rect 670 2358 674 2362
rect 726 2348 730 2352
rect 766 2338 770 2342
rect 662 2328 666 2332
rect 662 2318 666 2322
rect 694 2318 698 2322
rect 710 2318 714 2322
rect 694 2308 698 2312
rect 670 2278 674 2282
rect 574 2268 578 2272
rect 606 2268 610 2272
rect 654 2268 658 2272
rect 750 2308 754 2312
rect 742 2298 746 2302
rect 686 2268 690 2272
rect 734 2268 738 2272
rect 518 2258 522 2262
rect 510 2218 514 2222
rect 550 2198 554 2202
rect 518 2108 522 2112
rect 446 2088 450 2092
rect 470 2088 474 2092
rect 422 2078 426 2082
rect 430 2078 434 2082
rect 238 2058 242 2062
rect 246 2058 250 2062
rect 262 2058 266 2062
rect 318 2058 322 2062
rect 6 2048 10 2052
rect 54 2048 58 2052
rect 86 2048 90 2052
rect 6 2008 10 2012
rect 38 1988 42 1992
rect 70 1988 74 1992
rect 62 1968 66 1972
rect 78 1968 82 1972
rect 22 1958 26 1962
rect 54 1948 58 1952
rect 70 1948 74 1952
rect 142 1998 146 2002
rect 126 1978 130 1982
rect 222 1978 226 1982
rect 230 1968 234 1972
rect 238 1968 242 1972
rect 102 1958 106 1962
rect 134 1958 138 1962
rect 182 1958 186 1962
rect 206 1958 210 1962
rect 102 1948 106 1952
rect 86 1928 90 1932
rect 62 1898 66 1902
rect 30 1878 34 1882
rect 54 1878 58 1882
rect 158 1938 162 1942
rect 174 1938 178 1942
rect 166 1928 170 1932
rect 198 1928 202 1932
rect 190 1918 194 1922
rect 222 1938 226 1942
rect 230 1938 234 1942
rect 206 1898 210 1902
rect 110 1888 114 1892
rect 86 1878 90 1882
rect 102 1878 106 1882
rect 190 1878 194 1882
rect 30 1858 34 1862
rect 70 1858 74 1862
rect 6 1848 10 1852
rect 54 1848 58 1852
rect 86 1848 90 1852
rect 78 1828 82 1832
rect 30 1778 34 1782
rect 22 1758 26 1762
rect 6 1748 10 1752
rect 38 1688 42 1692
rect 6 1678 10 1682
rect 30 1658 34 1662
rect 394 2003 398 2007
rect 401 2003 405 2007
rect 350 1968 354 1972
rect 253 1948 257 1952
rect 334 1938 338 1942
rect 262 1918 266 1922
rect 366 1908 370 1912
rect 294 1888 298 1892
rect 398 1898 402 1902
rect 542 2108 546 2112
rect 670 2218 674 2222
rect 638 2208 642 2212
rect 614 2188 618 2192
rect 614 2178 618 2182
rect 614 2138 618 2142
rect 678 2138 682 2142
rect 630 2128 634 2132
rect 614 2108 618 2112
rect 654 2108 658 2112
rect 606 2078 610 2082
rect 646 2088 650 2092
rect 718 2258 722 2262
rect 886 2398 890 2402
rect 910 2398 914 2402
rect 862 2368 866 2372
rect 838 2348 842 2352
rect 822 2298 826 2302
rect 822 2278 826 2282
rect 766 2268 770 2272
rect 758 2258 762 2262
rect 814 2258 818 2262
rect 822 2258 826 2262
rect 838 2258 842 2262
rect 710 2248 714 2252
rect 822 2248 826 2252
rect 774 2228 778 2232
rect 878 2348 882 2352
rect 1014 2468 1018 2472
rect 1046 2468 1050 2472
rect 1054 2468 1058 2472
rect 1006 2338 1010 2342
rect 934 2328 938 2332
rect 982 2308 986 2312
rect 898 2303 902 2307
rect 905 2303 909 2307
rect 934 2298 938 2302
rect 902 2278 906 2282
rect 918 2268 922 2272
rect 878 2258 882 2262
rect 926 2258 930 2262
rect 878 2248 882 2252
rect 790 2238 794 2242
rect 846 2238 850 2242
rect 798 2228 802 2232
rect 862 2228 866 2232
rect 710 2188 714 2192
rect 702 2158 706 2162
rect 742 2178 746 2182
rect 814 2178 818 2182
rect 822 2178 826 2182
rect 846 2178 850 2182
rect 726 2168 730 2172
rect 734 2168 738 2172
rect 758 2168 762 2172
rect 798 2168 802 2172
rect 710 2138 714 2142
rect 686 2108 690 2112
rect 686 2098 690 2102
rect 726 2088 730 2092
rect 470 2068 474 2072
rect 502 2068 506 2072
rect 654 2068 658 2072
rect 478 2058 482 2062
rect 510 2058 514 2062
rect 526 2058 530 2062
rect 622 2058 626 2062
rect 446 1978 450 1982
rect 454 1938 458 1942
rect 430 1898 434 1902
rect 422 1888 426 1892
rect 382 1878 386 1882
rect 174 1848 178 1852
rect 278 1838 282 1842
rect 246 1788 250 1792
rect 262 1788 266 1792
rect 334 1768 338 1772
rect 158 1748 162 1752
rect 142 1738 146 1742
rect 158 1678 162 1682
rect 394 1803 398 1807
rect 401 1803 405 1807
rect 438 1858 442 1862
rect 462 1828 466 1832
rect 526 2048 530 2052
rect 630 2048 634 2052
rect 662 2048 666 2052
rect 486 2038 490 2042
rect 678 2028 682 2032
rect 630 2008 634 2012
rect 622 1998 626 2002
rect 662 1998 666 2002
rect 638 1978 642 1982
rect 654 1968 658 1972
rect 638 1958 642 1962
rect 694 1998 698 2002
rect 702 1988 706 1992
rect 686 1978 690 1982
rect 766 2148 770 2152
rect 758 2138 762 2142
rect 790 2138 794 2142
rect 750 2128 754 2132
rect 766 2128 770 2132
rect 814 2138 818 2142
rect 806 2108 810 2112
rect 798 2088 802 2092
rect 782 2068 786 2072
rect 758 2058 762 2062
rect 718 2048 722 2052
rect 774 2048 778 2052
rect 782 2048 786 2052
rect 686 1968 690 1972
rect 710 1968 714 1972
rect 542 1948 546 1952
rect 678 1948 682 1952
rect 526 1918 530 1922
rect 534 1878 538 1882
rect 550 1868 554 1872
rect 614 1938 618 1942
rect 638 1938 642 1942
rect 654 1938 658 1942
rect 686 1938 690 1942
rect 702 1938 706 1942
rect 710 1938 714 1942
rect 630 1908 634 1912
rect 654 1878 658 1882
rect 478 1858 482 1862
rect 470 1818 474 1822
rect 502 1798 506 1802
rect 438 1758 442 1762
rect 454 1758 458 1762
rect 270 1728 274 1732
rect 318 1718 322 1722
rect 214 1658 218 1662
rect 246 1658 250 1662
rect 230 1648 234 1652
rect 254 1648 258 1652
rect 142 1638 146 1642
rect 30 1588 34 1592
rect 6 1578 10 1582
rect 126 1578 130 1582
rect 22 1568 26 1572
rect 142 1568 146 1572
rect 238 1568 242 1572
rect 86 1558 90 1562
rect 70 1548 74 1552
rect 134 1548 138 1552
rect 6 1498 10 1502
rect 38 1498 42 1502
rect 30 1478 34 1482
rect 6 1468 10 1472
rect 6 1418 10 1422
rect 6 1378 10 1382
rect 22 1358 26 1362
rect 30 1348 34 1352
rect 62 1478 66 1482
rect 46 1468 50 1472
rect 142 1538 146 1542
rect 222 1538 226 1542
rect 166 1518 170 1522
rect 78 1498 82 1502
rect 78 1478 82 1482
rect 182 1478 186 1482
rect 78 1468 82 1472
rect 310 1638 314 1642
rect 382 1678 386 1682
rect 390 1678 394 1682
rect 342 1668 346 1672
rect 358 1668 362 1672
rect 382 1658 386 1662
rect 326 1638 330 1642
rect 318 1588 322 1592
rect 326 1578 330 1582
rect 310 1538 314 1542
rect 422 1668 426 1672
rect 470 1718 474 1722
rect 486 1718 490 1722
rect 614 1748 618 1752
rect 542 1738 546 1742
rect 542 1718 546 1722
rect 502 1678 506 1682
rect 430 1658 434 1662
rect 478 1658 482 1662
rect 398 1638 402 1642
rect 394 1603 398 1607
rect 401 1603 405 1607
rect 422 1598 426 1602
rect 366 1588 370 1592
rect 358 1498 362 1502
rect 398 1568 402 1572
rect 502 1638 506 1642
rect 526 1588 530 1592
rect 430 1548 434 1552
rect 382 1538 386 1542
rect 270 1478 274 1482
rect 302 1478 306 1482
rect 350 1478 354 1482
rect 46 1368 50 1372
rect 134 1398 138 1402
rect 94 1388 98 1392
rect 62 1378 66 1382
rect 102 1378 106 1382
rect 78 1368 82 1372
rect 182 1388 186 1392
rect 142 1378 146 1382
rect 126 1358 130 1362
rect 54 1348 58 1352
rect 110 1348 114 1352
rect 54 1338 58 1342
rect 102 1338 106 1342
rect 94 1268 98 1272
rect 110 1258 114 1262
rect 158 1258 162 1262
rect 54 1248 58 1252
rect 110 1248 114 1252
rect 126 1198 130 1202
rect 38 1168 42 1172
rect 94 1168 98 1172
rect 86 1158 90 1162
rect 62 1148 66 1152
rect 134 1148 138 1152
rect 126 1118 130 1122
rect 342 1398 346 1402
rect 254 1388 258 1392
rect 358 1388 362 1392
rect 350 1378 354 1382
rect 230 1358 234 1362
rect 302 1348 306 1352
rect 246 1328 250 1332
rect 214 1298 218 1302
rect 190 1258 194 1262
rect 158 1148 162 1152
rect 198 1148 202 1152
rect 150 1108 154 1112
rect 190 1098 194 1102
rect 6 1088 10 1092
rect 30 1078 34 1082
rect 158 1078 162 1082
rect 6 1068 10 1072
rect 142 1068 146 1072
rect 30 1058 34 1062
rect 6 1048 10 1052
rect 38 988 42 992
rect 6 978 10 982
rect 22 958 26 962
rect 158 948 162 952
rect 142 918 146 922
rect 142 888 146 892
rect 6 878 10 882
rect 30 858 34 862
rect 158 858 162 862
rect 22 848 26 852
rect 54 848 58 852
rect 46 838 50 842
rect 38 788 42 792
rect 6 778 10 782
rect 22 768 26 772
rect 158 748 162 752
rect 142 718 146 722
rect 166 708 170 712
rect 134 678 138 682
rect 6 648 10 652
rect 118 628 122 632
rect 134 628 138 632
rect 118 618 122 622
rect 14 538 18 542
rect 78 538 82 542
rect 6 448 10 452
rect 6 348 10 352
rect 62 478 66 482
rect 86 408 90 412
rect 94 388 98 392
rect 22 348 26 352
rect 14 338 18 342
rect 38 338 42 342
rect 6 148 10 152
rect 102 348 106 352
rect 150 608 154 612
rect 262 1288 266 1292
rect 478 1538 482 1542
rect 558 1708 562 1712
rect 654 1838 658 1842
rect 654 1778 658 1782
rect 710 1868 714 1872
rect 702 1858 706 1862
rect 742 2038 746 2042
rect 750 2038 754 2042
rect 742 1978 746 1982
rect 726 1968 730 1972
rect 766 1998 770 2002
rect 774 1978 778 1982
rect 758 1968 762 1972
rect 814 2058 818 2062
rect 870 2218 874 2222
rect 830 2168 834 2172
rect 838 2168 842 2172
rect 846 2148 850 2152
rect 838 2138 842 2142
rect 870 2138 874 2142
rect 958 2278 962 2282
rect 974 2278 978 2282
rect 1182 2638 1186 2642
rect 1150 2608 1154 2612
rect 1206 2648 1210 2652
rect 1126 2598 1130 2602
rect 1198 2598 1202 2602
rect 1110 2588 1114 2592
rect 1102 2558 1106 2562
rect 1094 2548 1098 2552
rect 1118 2548 1122 2552
rect 1366 2868 1370 2872
rect 1374 2848 1378 2852
rect 1350 2838 1354 2842
rect 1374 2838 1378 2842
rect 1270 2798 1274 2802
rect 1254 2768 1258 2772
rect 1246 2668 1250 2672
rect 1382 2808 1386 2812
rect 1414 2938 1418 2942
rect 1430 2938 1434 2942
rect 1558 2978 1562 2982
rect 1478 2968 1482 2972
rect 1534 2968 1538 2972
rect 1462 2958 1466 2962
rect 1534 2958 1538 2962
rect 1478 2948 1482 2952
rect 1422 2918 1426 2922
rect 1438 2918 1442 2922
rect 1398 2898 1402 2902
rect 1414 2888 1418 2892
rect 1430 2898 1434 2902
rect 1470 2938 1474 2942
rect 1486 2938 1490 2942
rect 1478 2928 1482 2932
rect 1494 2928 1498 2932
rect 1486 2908 1490 2912
rect 1454 2888 1458 2892
rect 1534 2938 1538 2942
rect 1542 2928 1546 2932
rect 1510 2918 1514 2922
rect 1558 2918 1562 2922
rect 1694 3098 1698 3102
rect 1930 3103 1934 3107
rect 1937 3103 1941 3107
rect 1902 3098 1906 3102
rect 1918 3098 1922 3102
rect 1894 3088 1898 3092
rect 1606 3058 1610 3062
rect 1582 2968 1586 2972
rect 1670 3058 1674 3062
rect 1838 3058 1842 3062
rect 1878 3058 1882 3062
rect 1638 2988 1642 2992
rect 1678 2948 1682 2952
rect 1574 2938 1578 2942
rect 1606 2938 1610 2942
rect 1622 2938 1626 2942
rect 1694 2938 1698 2942
rect 1582 2918 1586 2922
rect 1638 2928 1642 2932
rect 1598 2908 1602 2912
rect 1654 2908 1658 2912
rect 1702 2908 1706 2912
rect 1542 2888 1546 2892
rect 1638 2888 1642 2892
rect 1438 2878 1442 2882
rect 1494 2878 1498 2882
rect 1446 2858 1450 2862
rect 1462 2858 1466 2862
rect 1654 2858 1658 2862
rect 1418 2803 1422 2807
rect 1425 2803 1429 2807
rect 1390 2778 1394 2782
rect 1462 2848 1466 2852
rect 1502 2828 1506 2832
rect 1486 2808 1490 2812
rect 1350 2758 1354 2762
rect 1278 2748 1282 2752
rect 1262 2738 1266 2742
rect 1678 2848 1682 2852
rect 1670 2838 1674 2842
rect 1526 2788 1530 2792
rect 1542 2788 1546 2792
rect 1646 2768 1650 2772
rect 1782 2988 1786 2992
rect 1798 2998 1802 3002
rect 1790 2978 1794 2982
rect 1750 2928 1754 2932
rect 1718 2878 1722 2882
rect 1742 2878 1746 2882
rect 1814 2958 1818 2962
rect 1790 2878 1794 2882
rect 1878 2918 1882 2922
rect 1966 2928 1970 2932
rect 1894 2908 1898 2912
rect 1930 2903 1934 2907
rect 1937 2903 1941 2907
rect 1838 2898 1842 2902
rect 1886 2898 1890 2902
rect 1774 2868 1778 2872
rect 1814 2868 1818 2872
rect 1846 2868 1850 2872
rect 1950 2888 1954 2892
rect 1838 2858 1842 2862
rect 1934 2858 1938 2862
rect 1774 2848 1778 2852
rect 1750 2818 1754 2822
rect 1742 2808 1746 2812
rect 1686 2758 1690 2762
rect 1470 2748 1474 2752
rect 1494 2748 1498 2752
rect 1670 2748 1674 2752
rect 1694 2748 1698 2752
rect 1334 2728 1338 2732
rect 1262 2688 1266 2692
rect 1334 2678 1338 2682
rect 1430 2688 1434 2692
rect 1454 2668 1458 2672
rect 1350 2658 1354 2662
rect 1390 2658 1394 2662
rect 1262 2618 1266 2622
rect 1246 2588 1250 2592
rect 1326 2618 1330 2622
rect 1438 2618 1442 2622
rect 1278 2548 1282 2552
rect 1286 2548 1290 2552
rect 1142 2528 1146 2532
rect 1238 2528 1242 2532
rect 1078 2518 1082 2522
rect 1150 2498 1154 2502
rect 1238 2518 1242 2522
rect 1222 2488 1226 2492
rect 1086 2478 1090 2482
rect 1214 2478 1218 2482
rect 1070 2458 1074 2462
rect 1134 2458 1138 2462
rect 1062 2438 1066 2442
rect 1054 2338 1058 2342
rect 1030 2328 1034 2332
rect 1046 2308 1050 2312
rect 1206 2418 1210 2422
rect 1150 2408 1154 2412
rect 1126 2378 1130 2382
rect 1078 2368 1082 2372
rect 1094 2368 1098 2372
rect 1134 2368 1138 2372
rect 1078 2358 1082 2362
rect 1046 2288 1050 2292
rect 1054 2288 1058 2292
rect 1030 2278 1034 2282
rect 982 2268 986 2272
rect 950 2238 954 2242
rect 966 2228 970 2232
rect 942 2198 946 2202
rect 958 2168 962 2172
rect 966 2168 970 2172
rect 926 2148 930 2152
rect 958 2148 962 2152
rect 902 2138 906 2142
rect 918 2138 922 2142
rect 934 2138 938 2142
rect 878 2128 882 2132
rect 918 2128 922 2132
rect 886 2108 890 2112
rect 898 2103 902 2107
rect 905 2103 909 2107
rect 974 2118 978 2122
rect 862 2088 866 2092
rect 982 2088 986 2092
rect 942 2078 946 2082
rect 966 2078 970 2082
rect 854 2068 858 2072
rect 918 2068 922 2072
rect 806 2038 810 2042
rect 822 2038 826 2042
rect 806 2028 810 2032
rect 830 1998 834 2002
rect 814 1988 818 1992
rect 726 1878 730 1882
rect 742 1938 746 1942
rect 766 1918 770 1922
rect 790 1948 794 1952
rect 782 1918 786 1922
rect 734 1858 738 1862
rect 774 1878 778 1882
rect 878 2058 882 2062
rect 886 2038 890 2042
rect 862 1998 866 2002
rect 854 1988 858 1992
rect 878 1988 882 1992
rect 870 1978 874 1982
rect 822 1968 826 1972
rect 814 1948 818 1952
rect 838 1948 842 1952
rect 862 1948 866 1952
rect 870 1948 874 1952
rect 806 1898 810 1902
rect 950 2058 954 2062
rect 1006 2228 1010 2232
rect 1118 2358 1122 2362
rect 1102 2348 1106 2352
rect 1094 2328 1098 2332
rect 1086 2318 1090 2322
rect 1110 2308 1114 2312
rect 1038 2258 1042 2262
rect 1118 2258 1122 2262
rect 1022 2228 1026 2232
rect 1070 2228 1074 2232
rect 1094 2248 1098 2252
rect 1014 2168 1018 2172
rect 998 2158 1002 2162
rect 1014 2138 1018 2142
rect 998 2088 1002 2092
rect 990 2068 994 2072
rect 982 2058 986 2062
rect 1014 2058 1018 2062
rect 942 2018 946 2022
rect 934 1988 938 1992
rect 926 1978 930 1982
rect 910 1938 914 1942
rect 886 1908 890 1912
rect 898 1903 902 1907
rect 905 1903 909 1907
rect 886 1898 890 1902
rect 854 1878 858 1882
rect 862 1878 866 1882
rect 830 1868 834 1872
rect 862 1868 866 1872
rect 902 1878 906 1882
rect 886 1868 890 1872
rect 774 1858 778 1862
rect 798 1858 802 1862
rect 822 1858 826 1862
rect 846 1858 850 1862
rect 862 1858 866 1862
rect 878 1858 882 1862
rect 918 1858 922 1862
rect 758 1848 762 1852
rect 782 1848 786 1852
rect 702 1838 706 1842
rect 742 1838 746 1842
rect 742 1808 746 1812
rect 662 1768 666 1772
rect 694 1768 698 1772
rect 654 1748 658 1752
rect 638 1688 642 1692
rect 606 1678 610 1682
rect 590 1668 594 1672
rect 710 1738 714 1742
rect 694 1718 698 1722
rect 702 1708 706 1712
rect 774 1828 778 1832
rect 678 1688 682 1692
rect 742 1688 746 1692
rect 758 1688 762 1692
rect 718 1668 722 1672
rect 726 1668 730 1672
rect 662 1618 666 1622
rect 638 1598 642 1602
rect 582 1578 586 1582
rect 606 1578 610 1582
rect 630 1558 634 1562
rect 646 1578 650 1582
rect 718 1648 722 1652
rect 806 1818 810 1822
rect 814 1818 818 1822
rect 798 1808 802 1812
rect 790 1758 794 1762
rect 782 1728 786 1732
rect 758 1668 762 1672
rect 742 1648 746 1652
rect 750 1648 754 1652
rect 686 1638 690 1642
rect 702 1638 706 1642
rect 694 1578 698 1582
rect 694 1568 698 1572
rect 678 1558 682 1562
rect 614 1538 618 1542
rect 670 1538 674 1542
rect 694 1538 698 1542
rect 486 1518 490 1522
rect 518 1478 522 1482
rect 486 1468 490 1472
rect 510 1468 514 1472
rect 454 1438 458 1442
rect 438 1428 442 1432
rect 394 1403 398 1407
rect 401 1403 405 1407
rect 366 1358 370 1362
rect 374 1348 378 1352
rect 534 1468 538 1472
rect 502 1458 506 1462
rect 470 1378 474 1382
rect 502 1448 506 1452
rect 534 1438 538 1442
rect 534 1398 538 1402
rect 494 1348 498 1352
rect 518 1348 522 1352
rect 478 1318 482 1322
rect 462 1308 466 1312
rect 422 1298 426 1302
rect 398 1268 402 1272
rect 246 1258 250 1262
rect 366 1238 370 1242
rect 486 1268 490 1272
rect 518 1268 522 1272
rect 526 1268 530 1272
rect 430 1258 434 1262
rect 454 1258 458 1262
rect 502 1258 506 1262
rect 446 1248 450 1252
rect 478 1238 482 1242
rect 510 1238 514 1242
rect 534 1238 538 1242
rect 454 1218 458 1222
rect 414 1208 418 1212
rect 394 1203 398 1207
rect 401 1203 405 1207
rect 374 1178 378 1182
rect 406 1178 410 1182
rect 454 1178 458 1182
rect 358 1168 362 1172
rect 422 1168 426 1172
rect 430 1168 434 1172
rect 462 1168 466 1172
rect 502 1158 506 1162
rect 534 1158 538 1162
rect 374 1148 378 1152
rect 438 1148 442 1152
rect 222 1118 226 1122
rect 270 1118 274 1122
rect 254 1098 258 1102
rect 278 1088 282 1092
rect 534 1138 538 1142
rect 382 1118 386 1122
rect 366 1088 370 1092
rect 366 1078 370 1082
rect 246 1058 250 1062
rect 462 1128 466 1132
rect 430 1078 434 1082
rect 414 1068 418 1072
rect 422 1058 426 1062
rect 462 1058 466 1062
rect 350 1048 354 1052
rect 430 1048 434 1052
rect 430 1028 434 1032
rect 394 1003 398 1007
rect 401 1003 405 1007
rect 262 988 266 992
rect 302 988 306 992
rect 238 968 242 972
rect 286 968 290 972
rect 262 958 266 962
rect 390 978 394 982
rect 294 958 298 962
rect 494 1128 498 1132
rect 710 1588 714 1592
rect 726 1568 730 1572
rect 798 1688 802 1692
rect 758 1618 762 1622
rect 766 1598 770 1602
rect 766 1588 770 1592
rect 774 1568 778 1572
rect 742 1558 746 1562
rect 830 1828 834 1832
rect 830 1818 834 1822
rect 846 1778 850 1782
rect 894 1848 898 1852
rect 910 1828 914 1832
rect 870 1818 874 1822
rect 886 1768 890 1772
rect 950 1968 954 1972
rect 966 1948 970 1952
rect 990 2028 994 2032
rect 1006 2008 1010 2012
rect 982 1978 986 1982
rect 1038 2218 1042 2222
rect 1046 2208 1050 2212
rect 1030 2128 1034 2132
rect 1054 2128 1058 2132
rect 1038 2108 1042 2112
rect 1070 2168 1074 2172
rect 1110 2158 1114 2162
rect 1182 2398 1186 2402
rect 1158 2368 1162 2372
rect 1182 2368 1186 2372
rect 1158 2348 1162 2352
rect 1142 2338 1146 2342
rect 1270 2488 1274 2492
rect 1418 2603 1422 2607
rect 1425 2603 1429 2607
rect 1334 2558 1338 2562
rect 1390 2578 1394 2582
rect 1294 2528 1298 2532
rect 1430 2548 1434 2552
rect 1486 2708 1490 2712
rect 1478 2678 1482 2682
rect 1478 2668 1482 2672
rect 1470 2618 1474 2622
rect 1406 2488 1410 2492
rect 1462 2488 1466 2492
rect 1286 2478 1290 2482
rect 1438 2478 1442 2482
rect 1278 2468 1282 2472
rect 1366 2468 1370 2472
rect 1430 2468 1434 2472
rect 1614 2728 1618 2732
rect 1558 2698 1562 2702
rect 1582 2698 1586 2702
rect 1526 2678 1530 2682
rect 1542 2668 1546 2672
rect 1542 2648 1546 2652
rect 1582 2608 1586 2612
rect 1518 2558 1522 2562
rect 1502 2528 1506 2532
rect 1518 2508 1522 2512
rect 1518 2468 1522 2472
rect 1326 2458 1330 2462
rect 1358 2458 1362 2462
rect 1374 2458 1378 2462
rect 1470 2458 1474 2462
rect 1270 2438 1274 2442
rect 1302 2438 1306 2442
rect 1230 2408 1234 2412
rect 1342 2448 1346 2452
rect 1374 2448 1378 2452
rect 1366 2438 1370 2442
rect 1318 2428 1322 2432
rect 1310 2368 1314 2372
rect 1334 2418 1338 2422
rect 1318 2348 1322 2352
rect 1206 2338 1210 2342
rect 1174 2318 1178 2322
rect 1270 2338 1274 2342
rect 1318 2338 1322 2342
rect 1254 2328 1258 2332
rect 1318 2308 1322 2312
rect 1214 2298 1218 2302
rect 1246 2298 1250 2302
rect 1350 2398 1354 2402
rect 1342 2358 1346 2362
rect 1342 2348 1346 2352
rect 1318 2278 1322 2282
rect 1310 2268 1314 2272
rect 1190 2258 1194 2262
rect 1174 2208 1178 2212
rect 1158 2188 1162 2192
rect 1078 2138 1082 2142
rect 1094 2138 1098 2142
rect 1118 2138 1122 2142
rect 1070 2128 1074 2132
rect 1054 2098 1058 2102
rect 1062 2098 1066 2102
rect 1142 2118 1146 2122
rect 1078 2108 1082 2112
rect 1118 2108 1122 2112
rect 1062 2088 1066 2092
rect 1046 2058 1050 2062
rect 1070 2058 1074 2062
rect 1102 2058 1106 2062
rect 1030 2028 1034 2032
rect 1030 2008 1034 2012
rect 1038 1998 1042 2002
rect 1054 1998 1058 2002
rect 1014 1968 1018 1972
rect 998 1958 1002 1962
rect 1030 1948 1034 1952
rect 982 1938 986 1942
rect 998 1938 1002 1942
rect 1022 1938 1026 1942
rect 974 1908 978 1912
rect 974 1898 978 1902
rect 1014 1888 1018 1892
rect 1006 1878 1010 1882
rect 958 1868 962 1872
rect 966 1858 970 1862
rect 982 1858 986 1862
rect 958 1808 962 1812
rect 934 1768 938 1772
rect 950 1768 954 1772
rect 910 1748 914 1752
rect 926 1748 930 1752
rect 830 1738 834 1742
rect 870 1738 874 1742
rect 814 1698 818 1702
rect 838 1728 842 1732
rect 918 1728 922 1732
rect 862 1718 866 1722
rect 846 1698 850 1702
rect 822 1658 826 1662
rect 790 1648 794 1652
rect 814 1568 818 1572
rect 766 1548 770 1552
rect 814 1548 818 1552
rect 742 1528 746 1532
rect 782 1498 786 1502
rect 566 1478 570 1482
rect 670 1478 674 1482
rect 718 1478 722 1482
rect 630 1468 634 1472
rect 646 1468 650 1472
rect 726 1468 730 1472
rect 758 1468 762 1472
rect 798 1468 802 1472
rect 606 1458 610 1462
rect 638 1458 642 1462
rect 654 1458 658 1462
rect 750 1458 754 1462
rect 790 1458 794 1462
rect 566 1448 570 1452
rect 558 1438 562 1442
rect 590 1438 594 1442
rect 550 1428 554 1432
rect 598 1428 602 1432
rect 646 1428 650 1432
rect 574 1398 578 1402
rect 606 1398 610 1402
rect 574 1328 578 1332
rect 590 1288 594 1292
rect 550 1278 554 1282
rect 590 1278 594 1282
rect 566 1258 570 1262
rect 574 1238 578 1242
rect 558 1208 562 1212
rect 558 1198 562 1202
rect 550 1178 554 1182
rect 678 1438 682 1442
rect 694 1438 698 1442
rect 798 1438 802 1442
rect 686 1428 690 1432
rect 686 1418 690 1422
rect 686 1388 690 1392
rect 670 1368 674 1372
rect 678 1338 682 1342
rect 662 1288 666 1292
rect 622 1268 626 1272
rect 630 1268 634 1272
rect 654 1268 658 1272
rect 670 1268 674 1272
rect 598 1258 602 1262
rect 614 1258 618 1262
rect 630 1248 634 1252
rect 582 1228 586 1232
rect 614 1208 618 1212
rect 590 1178 594 1182
rect 566 1168 570 1172
rect 582 1168 586 1172
rect 686 1298 690 1302
rect 918 1708 922 1712
rect 898 1703 902 1707
rect 905 1703 909 1707
rect 870 1678 874 1682
rect 894 1678 898 1682
rect 878 1658 882 1662
rect 942 1738 946 1742
rect 950 1728 954 1732
rect 934 1718 938 1722
rect 1110 2038 1114 2042
rect 1086 2028 1090 2032
rect 1078 1988 1082 1992
rect 1070 1968 1074 1972
rect 1054 1948 1058 1952
rect 1070 1948 1074 1952
rect 1102 1978 1106 1982
rect 1086 1938 1090 1942
rect 1038 1878 1042 1882
rect 1134 2088 1138 2092
rect 1126 2048 1130 2052
rect 1142 2038 1146 2042
rect 1126 2028 1130 2032
rect 1158 2048 1162 2052
rect 1150 2018 1154 2022
rect 1126 2008 1130 2012
rect 1158 2008 1162 2012
rect 1102 1908 1106 1912
rect 1038 1858 1042 1862
rect 1054 1858 1058 1862
rect 1078 1858 1082 1862
rect 1094 1858 1098 1862
rect 974 1828 978 1832
rect 998 1828 1002 1832
rect 1030 1828 1034 1832
rect 1006 1758 1010 1762
rect 990 1738 994 1742
rect 990 1728 994 1732
rect 942 1688 946 1692
rect 966 1688 970 1692
rect 982 1688 986 1692
rect 902 1658 906 1662
rect 918 1658 922 1662
rect 926 1658 930 1662
rect 950 1648 954 1652
rect 838 1638 842 1642
rect 878 1628 882 1632
rect 830 1618 834 1622
rect 886 1598 890 1602
rect 846 1588 850 1592
rect 838 1578 842 1582
rect 814 1468 818 1472
rect 822 1428 826 1432
rect 878 1578 882 1582
rect 886 1578 890 1582
rect 870 1548 874 1552
rect 846 1498 850 1502
rect 854 1498 858 1502
rect 838 1478 842 1482
rect 982 1668 986 1672
rect 942 1638 946 1642
rect 958 1638 962 1642
rect 974 1638 978 1642
rect 910 1588 914 1592
rect 958 1578 962 1582
rect 942 1568 946 1572
rect 894 1558 898 1562
rect 982 1568 986 1572
rect 894 1548 898 1552
rect 966 1548 970 1552
rect 974 1548 978 1552
rect 870 1528 874 1532
rect 870 1518 874 1522
rect 870 1508 874 1512
rect 898 1503 902 1507
rect 905 1503 909 1507
rect 878 1468 882 1472
rect 886 1468 890 1472
rect 902 1468 906 1472
rect 878 1448 882 1452
rect 926 1488 930 1492
rect 918 1438 922 1442
rect 846 1428 850 1432
rect 870 1428 874 1432
rect 806 1418 810 1422
rect 702 1348 706 1352
rect 758 1408 762 1412
rect 782 1408 786 1412
rect 766 1398 770 1402
rect 750 1378 754 1382
rect 806 1398 810 1402
rect 798 1378 802 1382
rect 734 1358 738 1362
rect 862 1408 866 1412
rect 846 1378 850 1382
rect 854 1368 858 1372
rect 846 1358 850 1362
rect 862 1358 866 1362
rect 790 1348 794 1352
rect 806 1348 810 1352
rect 830 1348 834 1352
rect 838 1348 842 1352
rect 710 1338 714 1342
rect 750 1338 754 1342
rect 718 1298 722 1302
rect 702 1278 706 1282
rect 678 1258 682 1262
rect 710 1258 714 1262
rect 654 1248 658 1252
rect 662 1248 666 1252
rect 710 1248 714 1252
rect 638 1218 642 1222
rect 646 1178 650 1182
rect 638 1158 642 1162
rect 606 1128 610 1132
rect 542 1118 546 1122
rect 574 1118 578 1122
rect 550 1098 554 1102
rect 534 1088 538 1092
rect 518 1078 522 1082
rect 518 1048 522 1052
rect 614 1108 618 1112
rect 606 1068 610 1072
rect 534 1008 538 1012
rect 478 978 482 982
rect 478 968 482 972
rect 582 948 586 952
rect 438 938 442 942
rect 510 938 514 942
rect 526 938 530 942
rect 622 938 626 942
rect 374 918 378 922
rect 262 878 266 882
rect 454 878 458 882
rect 238 868 242 872
rect 302 868 306 872
rect 214 728 218 732
rect 254 858 258 862
rect 238 848 242 852
rect 230 778 234 782
rect 326 838 330 842
rect 318 768 322 772
rect 270 738 274 742
rect 286 738 290 742
rect 222 708 226 712
rect 230 688 234 692
rect 302 708 306 712
rect 366 838 370 842
rect 394 803 398 807
rect 401 803 405 807
rect 390 778 394 782
rect 422 778 426 782
rect 342 738 346 742
rect 366 738 370 742
rect 310 698 314 702
rect 566 898 570 902
rect 550 868 554 872
rect 438 708 442 712
rect 550 848 554 852
rect 558 848 562 852
rect 534 808 538 812
rect 526 748 530 752
rect 622 888 626 892
rect 646 1128 650 1132
rect 742 1328 746 1332
rect 742 1318 746 1322
rect 758 1318 762 1322
rect 750 1308 754 1312
rect 766 1308 770 1312
rect 838 1328 842 1332
rect 822 1308 826 1312
rect 790 1298 794 1302
rect 862 1338 866 1342
rect 854 1298 858 1302
rect 774 1288 778 1292
rect 822 1288 826 1292
rect 830 1268 834 1272
rect 734 1258 738 1262
rect 726 1208 730 1212
rect 694 1198 698 1202
rect 702 1158 706 1162
rect 686 1148 690 1152
rect 702 1148 706 1152
rect 718 1148 722 1152
rect 670 1128 674 1132
rect 678 1118 682 1122
rect 670 1098 674 1102
rect 654 1078 658 1082
rect 662 1078 666 1082
rect 638 1068 642 1072
rect 654 1068 658 1072
rect 646 1058 650 1062
rect 638 938 642 942
rect 718 1118 722 1122
rect 742 1228 746 1232
rect 766 1198 770 1202
rect 750 1168 754 1172
rect 774 1168 778 1172
rect 766 1148 770 1152
rect 750 1128 754 1132
rect 734 1108 738 1112
rect 726 1068 730 1072
rect 734 1068 738 1072
rect 766 1068 770 1072
rect 742 1058 746 1062
rect 662 1048 666 1052
rect 678 1048 682 1052
rect 702 1048 706 1052
rect 718 1048 722 1052
rect 774 1048 778 1052
rect 662 1038 666 1042
rect 670 1018 674 1022
rect 662 938 666 942
rect 654 928 658 932
rect 582 808 586 812
rect 614 808 618 812
rect 566 738 570 742
rect 558 728 562 732
rect 478 708 482 712
rect 422 698 426 702
rect 438 698 442 702
rect 454 698 458 702
rect 470 698 474 702
rect 382 678 386 682
rect 198 668 202 672
rect 326 668 330 672
rect 190 658 194 662
rect 230 658 234 662
rect 150 558 154 562
rect 190 548 194 552
rect 174 538 178 542
rect 142 528 146 532
rect 190 528 194 532
rect 182 468 186 472
rect 118 318 122 322
rect 142 318 146 322
rect 94 278 98 282
rect 110 258 114 262
rect 38 188 42 192
rect 54 188 58 192
rect 78 188 82 192
rect 278 618 282 622
rect 394 603 398 607
rect 401 603 405 607
rect 278 578 282 582
rect 406 568 410 572
rect 470 678 474 682
rect 438 558 442 562
rect 430 548 434 552
rect 422 538 426 542
rect 398 528 402 532
rect 294 518 298 522
rect 286 488 290 492
rect 230 458 234 462
rect 270 458 274 462
rect 214 388 218 392
rect 302 358 306 362
rect 406 438 410 442
rect 374 428 378 432
rect 394 403 398 407
rect 401 403 405 407
rect 390 368 394 372
rect 262 348 266 352
rect 278 348 282 352
rect 326 348 330 352
rect 334 348 338 352
rect 206 328 210 332
rect 358 308 362 312
rect 190 298 194 302
rect 262 288 266 292
rect 150 258 154 262
rect 190 258 194 262
rect 406 298 410 302
rect 374 288 378 292
rect 534 688 538 692
rect 510 668 514 672
rect 542 558 546 562
rect 598 758 602 762
rect 702 1038 706 1042
rect 726 1038 730 1042
rect 750 1038 754 1042
rect 710 1018 714 1022
rect 838 1258 842 1262
rect 822 1248 826 1252
rect 846 1248 850 1252
rect 838 1238 842 1242
rect 798 1188 802 1192
rect 790 1158 794 1162
rect 814 1168 818 1172
rect 894 1408 898 1412
rect 902 1358 906 1362
rect 918 1358 922 1362
rect 918 1348 922 1352
rect 942 1368 946 1372
rect 894 1338 898 1342
rect 934 1318 938 1322
rect 898 1303 902 1307
rect 905 1303 909 1307
rect 886 1288 890 1292
rect 942 1288 946 1292
rect 966 1528 970 1532
rect 958 1508 962 1512
rect 1022 1758 1026 1762
rect 1062 1818 1066 1822
rect 1078 1818 1082 1822
rect 1062 1768 1066 1772
rect 1038 1738 1042 1742
rect 1046 1738 1050 1742
rect 1054 1728 1058 1732
rect 1014 1718 1018 1722
rect 998 1658 1002 1662
rect 1006 1628 1010 1632
rect 998 1598 1002 1602
rect 990 1508 994 1512
rect 974 1468 978 1472
rect 990 1458 994 1462
rect 982 1448 986 1452
rect 966 1438 970 1442
rect 966 1308 970 1312
rect 974 1298 978 1302
rect 878 1268 882 1272
rect 886 1268 890 1272
rect 934 1268 938 1272
rect 854 1208 858 1212
rect 950 1258 954 1262
rect 910 1228 914 1232
rect 918 1218 922 1222
rect 918 1178 922 1182
rect 926 1178 930 1182
rect 854 1158 858 1162
rect 950 1158 954 1162
rect 1006 1548 1010 1552
rect 1022 1648 1026 1652
rect 1022 1598 1026 1602
rect 1038 1718 1042 1722
rect 1118 1908 1122 1912
rect 1110 1878 1114 1882
rect 1110 1858 1114 1862
rect 1102 1818 1106 1822
rect 1358 2338 1362 2342
rect 1326 2238 1330 2242
rect 1318 2228 1322 2232
rect 1278 2218 1282 2222
rect 1286 2198 1290 2202
rect 1182 2078 1186 2082
rect 1230 2138 1234 2142
rect 1246 2128 1250 2132
rect 1198 2098 1202 2102
rect 1230 2098 1234 2102
rect 1206 2088 1210 2092
rect 1190 2058 1194 2062
rect 1318 2158 1322 2162
rect 1310 2138 1314 2142
rect 1270 2078 1274 2082
rect 1214 2058 1218 2062
rect 1270 2058 1274 2062
rect 1190 2048 1194 2052
rect 1182 1978 1186 1982
rect 1134 1958 1138 1962
rect 1158 1958 1162 1962
rect 1166 1948 1170 1952
rect 1150 1938 1154 1942
rect 1166 1938 1170 1942
rect 1158 1888 1162 1892
rect 1174 1868 1178 1872
rect 1142 1858 1146 1862
rect 1230 2018 1234 2022
rect 1262 1988 1266 1992
rect 1254 1968 1258 1972
rect 1262 1968 1266 1972
rect 1214 1948 1218 1952
rect 1238 1938 1242 1942
rect 1198 1928 1202 1932
rect 1238 1918 1242 1922
rect 1222 1908 1226 1912
rect 1214 1878 1218 1882
rect 1222 1858 1226 1862
rect 1134 1838 1138 1842
rect 1134 1818 1138 1822
rect 1166 1828 1170 1832
rect 1150 1788 1154 1792
rect 1110 1768 1114 1772
rect 1126 1768 1130 1772
rect 1142 1758 1146 1762
rect 1150 1758 1154 1762
rect 1078 1728 1082 1732
rect 1070 1718 1074 1722
rect 1118 1738 1122 1742
rect 1102 1708 1106 1712
rect 1142 1708 1146 1712
rect 1094 1678 1098 1682
rect 1262 1958 1266 1962
rect 1254 1878 1258 1882
rect 1222 1838 1226 1842
rect 1222 1808 1226 1812
rect 1182 1788 1186 1792
rect 1230 1788 1234 1792
rect 1230 1778 1234 1782
rect 1182 1768 1186 1772
rect 1302 1978 1306 1982
rect 1318 1978 1322 1982
rect 1310 1968 1314 1972
rect 1278 1948 1282 1952
rect 1334 2128 1338 2132
rect 1382 2418 1386 2422
rect 1454 2418 1458 2422
rect 1438 2408 1442 2412
rect 1418 2403 1422 2407
rect 1425 2403 1429 2407
rect 1398 2388 1402 2392
rect 1462 2398 1466 2402
rect 1454 2358 1458 2362
rect 1390 2348 1394 2352
rect 1486 2448 1490 2452
rect 1502 2448 1506 2452
rect 1518 2438 1522 2442
rect 1494 2428 1498 2432
rect 1502 2428 1506 2432
rect 1574 2538 1578 2542
rect 1630 2688 1634 2692
rect 1686 2688 1690 2692
rect 1646 2678 1650 2682
rect 1654 2668 1658 2672
rect 1846 2848 1850 2852
rect 1790 2838 1794 2842
rect 1782 2828 1786 2832
rect 1774 2798 1778 2802
rect 1750 2748 1754 2752
rect 1814 2728 1818 2732
rect 1798 2718 1802 2722
rect 1734 2678 1738 2682
rect 1630 2648 1634 2652
rect 1654 2608 1658 2612
rect 1862 2828 1866 2832
rect 1878 2808 1882 2812
rect 1870 2778 1874 2782
rect 2062 3038 2066 3042
rect 2030 2988 2034 2992
rect 2046 2988 2050 2992
rect 2038 2938 2042 2942
rect 2038 2908 2042 2912
rect 2030 2898 2034 2902
rect 2142 3098 2146 3102
rect 2174 3098 2178 3102
rect 2086 3058 2090 3062
rect 2126 3058 2130 3062
rect 2086 3018 2090 3022
rect 2078 2988 2082 2992
rect 2174 3008 2178 3012
rect 2190 2988 2194 2992
rect 2086 2948 2090 2952
rect 2182 2948 2186 2952
rect 2062 2938 2066 2942
rect 2054 2898 2058 2902
rect 2166 2918 2170 2922
rect 2174 2908 2178 2912
rect 2158 2858 2162 2862
rect 2070 2828 2074 2832
rect 1998 2818 2002 2822
rect 1886 2778 1890 2782
rect 1886 2768 1890 2772
rect 1990 2758 1994 2762
rect 2094 2758 2098 2762
rect 2094 2748 2098 2752
rect 2214 2768 2218 2772
rect 2134 2758 2138 2762
rect 2198 2758 2202 2762
rect 2158 2748 2162 2752
rect 2006 2728 2010 2732
rect 2054 2728 2058 2732
rect 2102 2728 2106 2732
rect 1910 2718 1914 2722
rect 1930 2703 1934 2707
rect 1937 2703 1941 2707
rect 1926 2678 1930 2682
rect 1910 2668 1914 2672
rect 2046 2668 2050 2672
rect 1886 2658 1890 2662
rect 1902 2658 1906 2662
rect 2046 2658 2050 2662
rect 1854 2638 1858 2642
rect 1806 2618 1810 2622
rect 1766 2608 1770 2612
rect 1782 2578 1786 2582
rect 1750 2568 1754 2572
rect 1614 2548 1618 2552
rect 1758 2548 1762 2552
rect 1774 2548 1778 2552
rect 1822 2608 1826 2612
rect 1830 2558 1834 2562
rect 1854 2588 1858 2592
rect 1894 2578 1898 2582
rect 1894 2558 1898 2562
rect 1942 2558 1946 2562
rect 1838 2548 1842 2552
rect 1878 2548 1882 2552
rect 1782 2538 1786 2542
rect 1598 2528 1602 2532
rect 1558 2518 1562 2522
rect 1766 2528 1770 2532
rect 1670 2518 1674 2522
rect 1630 2508 1634 2512
rect 1654 2508 1658 2512
rect 1670 2488 1674 2492
rect 1734 2488 1738 2492
rect 1790 2498 1794 2502
rect 1798 2498 1802 2502
rect 1678 2478 1682 2482
rect 1694 2478 1698 2482
rect 1702 2478 1706 2482
rect 1718 2478 1722 2482
rect 1598 2468 1602 2472
rect 1630 2468 1634 2472
rect 1646 2468 1650 2472
rect 1654 2458 1658 2462
rect 1542 2448 1546 2452
rect 1582 2448 1586 2452
rect 1614 2448 1618 2452
rect 1566 2438 1570 2442
rect 1582 2438 1586 2442
rect 1630 2438 1634 2442
rect 1646 2438 1650 2442
rect 1550 2428 1554 2432
rect 1638 2428 1642 2432
rect 1662 2428 1666 2432
rect 1582 2418 1586 2422
rect 1526 2408 1530 2412
rect 1478 2388 1482 2392
rect 1526 2388 1530 2392
rect 1494 2348 1498 2352
rect 1534 2348 1538 2352
rect 1382 2338 1386 2342
rect 1406 2338 1410 2342
rect 1502 2338 1506 2342
rect 1542 2338 1546 2342
rect 1390 2298 1394 2302
rect 1382 2208 1386 2212
rect 1390 2188 1394 2192
rect 1382 2168 1386 2172
rect 1342 2078 1346 2082
rect 1366 2138 1370 2142
rect 1358 2128 1362 2132
rect 1398 2178 1402 2182
rect 1478 2328 1482 2332
rect 1454 2318 1458 2322
rect 1446 2298 1450 2302
rect 1494 2308 1498 2312
rect 1510 2288 1514 2292
rect 1438 2278 1442 2282
rect 1418 2203 1422 2207
rect 1425 2203 1429 2207
rect 1430 2158 1434 2162
rect 1414 2128 1418 2132
rect 1518 2258 1522 2262
rect 1446 2218 1450 2222
rect 1406 2108 1410 2112
rect 1438 2108 1442 2112
rect 1358 2048 1362 2052
rect 1350 2018 1354 2022
rect 1342 1978 1346 1982
rect 1814 2508 1818 2512
rect 1806 2488 1810 2492
rect 1710 2468 1714 2472
rect 1750 2468 1754 2472
rect 1870 2518 1874 2522
rect 1870 2478 1874 2482
rect 1878 2478 1882 2482
rect 1830 2458 1834 2462
rect 1862 2458 1866 2462
rect 1806 2448 1810 2452
rect 1742 2438 1746 2442
rect 1774 2438 1778 2442
rect 1710 2428 1714 2432
rect 1742 2428 1746 2432
rect 1686 2408 1690 2412
rect 1678 2398 1682 2402
rect 1654 2358 1658 2362
rect 1662 2348 1666 2352
rect 1750 2408 1754 2412
rect 1734 2388 1738 2392
rect 1686 2358 1690 2362
rect 1710 2358 1714 2362
rect 1718 2348 1722 2352
rect 1758 2398 1762 2402
rect 1798 2428 1802 2432
rect 1822 2428 1826 2432
rect 1750 2368 1754 2372
rect 1774 2368 1778 2372
rect 1806 2378 1810 2382
rect 1806 2368 1810 2372
rect 1750 2358 1754 2362
rect 1790 2358 1794 2362
rect 1814 2358 1818 2362
rect 1758 2348 1762 2352
rect 1774 2348 1778 2352
rect 1798 2348 1802 2352
rect 1654 2338 1658 2342
rect 1670 2338 1674 2342
rect 1694 2338 1698 2342
rect 1718 2338 1722 2342
rect 1606 2328 1610 2332
rect 1646 2328 1650 2332
rect 1622 2318 1626 2322
rect 1598 2288 1602 2292
rect 1590 2278 1594 2282
rect 1606 2278 1610 2282
rect 1638 2278 1642 2282
rect 1606 2258 1610 2262
rect 1550 2248 1554 2252
rect 1566 2238 1570 2242
rect 1630 2248 1634 2252
rect 1606 2228 1610 2232
rect 1518 2218 1522 2222
rect 1542 2218 1546 2222
rect 1534 2208 1538 2212
rect 1606 2208 1610 2212
rect 1494 2198 1498 2202
rect 1510 2198 1514 2202
rect 1526 2138 1530 2142
rect 1486 2108 1490 2112
rect 1494 2098 1498 2102
rect 1406 2078 1410 2082
rect 1382 2068 1386 2072
rect 1470 2068 1474 2072
rect 1462 2058 1466 2062
rect 1502 2058 1506 2062
rect 1382 2038 1386 2042
rect 1398 2028 1402 2032
rect 1438 2028 1442 2032
rect 1390 1998 1394 2002
rect 1382 1988 1386 1992
rect 1374 1958 1378 1962
rect 1326 1948 1330 1952
rect 1278 1938 1282 1942
rect 1358 1938 1362 1942
rect 1342 1928 1346 1932
rect 1350 1928 1354 1932
rect 1310 1908 1314 1912
rect 1294 1878 1298 1882
rect 1334 1878 1338 1882
rect 1390 1938 1394 1942
rect 1366 1888 1370 1892
rect 1326 1868 1330 1872
rect 1270 1858 1274 1862
rect 1278 1858 1282 1862
rect 1302 1858 1306 1862
rect 1358 1858 1362 1862
rect 1254 1838 1258 1842
rect 1262 1828 1266 1832
rect 1262 1788 1266 1792
rect 1270 1788 1274 1792
rect 1198 1758 1202 1762
rect 1246 1758 1250 1762
rect 1174 1738 1178 1742
rect 1198 1738 1202 1742
rect 1286 1778 1290 1782
rect 1270 1748 1274 1752
rect 1366 1838 1370 1842
rect 1334 1828 1338 1832
rect 1350 1828 1354 1832
rect 1358 1828 1362 1832
rect 1326 1778 1330 1782
rect 1302 1768 1306 1772
rect 1302 1758 1306 1762
rect 1294 1748 1298 1752
rect 1342 1748 1346 1752
rect 1214 1738 1218 1742
rect 1246 1738 1250 1742
rect 1206 1728 1210 1732
rect 1174 1678 1178 1682
rect 1038 1668 1042 1672
rect 1198 1668 1202 1672
rect 1046 1658 1050 1662
rect 1086 1648 1090 1652
rect 1230 1728 1234 1732
rect 1262 1728 1266 1732
rect 1390 1908 1394 1912
rect 1382 1828 1386 1832
rect 1390 1828 1394 1832
rect 1374 1818 1378 1822
rect 1374 1798 1378 1802
rect 1418 2003 1422 2007
rect 1425 2003 1429 2007
rect 1462 2008 1466 2012
rect 1438 1958 1442 1962
rect 1470 1978 1474 1982
rect 1438 1938 1442 1942
rect 1462 1928 1466 1932
rect 1406 1908 1410 1912
rect 1446 1908 1450 1912
rect 1486 1928 1490 1932
rect 1478 1908 1482 1912
rect 1478 1898 1482 1902
rect 1406 1878 1410 1882
rect 1454 1878 1458 1882
rect 1470 1878 1474 1882
rect 1462 1848 1466 1852
rect 1422 1838 1426 1842
rect 1446 1838 1450 1842
rect 1406 1808 1410 1812
rect 1438 1808 1442 1812
rect 1418 1803 1422 1807
rect 1425 1803 1429 1807
rect 1534 2098 1538 2102
rect 1526 2078 1530 2082
rect 1510 1898 1514 1902
rect 1566 2078 1570 2082
rect 1598 2078 1602 2082
rect 1662 2278 1666 2282
rect 1694 2308 1698 2312
rect 1678 2298 1682 2302
rect 1710 2298 1714 2302
rect 1758 2328 1762 2332
rect 1766 2328 1770 2332
rect 1774 2308 1778 2312
rect 1750 2298 1754 2302
rect 1702 2278 1706 2282
rect 1726 2278 1730 2282
rect 1734 2268 1738 2272
rect 1670 2258 1674 2262
rect 1758 2258 1762 2262
rect 1654 2198 1658 2202
rect 1630 2188 1634 2192
rect 1614 2148 1618 2152
rect 1694 2248 1698 2252
rect 1782 2248 1786 2252
rect 1686 2238 1690 2242
rect 1758 2228 1762 2232
rect 1782 2228 1786 2232
rect 1694 2208 1698 2212
rect 1662 2188 1666 2192
rect 1686 2168 1690 2172
rect 1742 2168 1746 2172
rect 1838 2418 1842 2422
rect 1830 2398 1834 2402
rect 1830 2358 1834 2362
rect 1814 2328 1818 2332
rect 1806 2278 1810 2282
rect 1814 2238 1818 2242
rect 1886 2468 1890 2472
rect 1910 2538 1914 2542
rect 1990 2598 1994 2602
rect 2006 2538 2010 2542
rect 2022 2538 2026 2542
rect 1950 2518 1954 2522
rect 1930 2503 1934 2507
rect 1937 2503 1941 2507
rect 1918 2498 1922 2502
rect 1934 2468 1938 2472
rect 1958 2498 1962 2502
rect 2118 2738 2122 2742
rect 2142 2728 2146 2732
rect 2110 2688 2114 2692
rect 2142 2668 2146 2672
rect 2166 2728 2170 2732
rect 2230 2748 2234 2752
rect 2222 2738 2226 2742
rect 2230 2708 2234 2712
rect 2166 2668 2170 2672
rect 2406 3098 2410 3102
rect 2486 3098 2490 3102
rect 2510 3088 2514 3092
rect 2406 3068 2410 3072
rect 2318 3018 2322 3022
rect 2438 3018 2442 3022
rect 2270 2968 2274 2972
rect 2254 2958 2258 2962
rect 2278 2958 2282 2962
rect 2294 2958 2298 2962
rect 2254 2788 2258 2792
rect 2286 2878 2290 2882
rect 2302 2928 2306 2932
rect 2442 3003 2446 3007
rect 2449 3003 2453 3007
rect 2342 2948 2346 2952
rect 2398 2948 2402 2952
rect 2470 2948 2474 2952
rect 2478 2948 2482 2952
rect 2326 2898 2330 2902
rect 2334 2878 2338 2882
rect 2310 2868 2314 2872
rect 2294 2848 2298 2852
rect 2414 2908 2418 2912
rect 2422 2898 2426 2902
rect 2350 2828 2354 2832
rect 2494 2928 2498 2932
rect 2486 2838 2490 2842
rect 2358 2818 2362 2822
rect 2382 2818 2386 2822
rect 2438 2818 2442 2822
rect 2342 2798 2346 2802
rect 2262 2768 2266 2772
rect 2302 2758 2306 2762
rect 2462 2808 2466 2812
rect 2442 2803 2446 2807
rect 2449 2803 2453 2807
rect 2414 2798 2418 2802
rect 2318 2738 2322 2742
rect 2270 2718 2274 2722
rect 2254 2678 2258 2682
rect 2478 2768 2482 2772
rect 2438 2748 2442 2752
rect 2422 2718 2426 2722
rect 2398 2708 2402 2712
rect 2406 2708 2410 2712
rect 2358 2698 2362 2702
rect 2318 2688 2322 2692
rect 2366 2678 2370 2682
rect 2382 2678 2386 2682
rect 2398 2678 2402 2682
rect 2358 2668 2362 2672
rect 2134 2658 2138 2662
rect 2150 2658 2154 2662
rect 2190 2658 2194 2662
rect 2230 2658 2234 2662
rect 2270 2658 2274 2662
rect 2302 2658 2306 2662
rect 2318 2658 2322 2662
rect 2334 2658 2338 2662
rect 2350 2658 2354 2662
rect 2142 2638 2146 2642
rect 2158 2638 2162 2642
rect 2190 2638 2194 2642
rect 2174 2618 2178 2622
rect 2166 2598 2170 2602
rect 2078 2558 2082 2562
rect 2094 2558 2098 2562
rect 2110 2558 2114 2562
rect 2174 2558 2178 2562
rect 2078 2548 2082 2552
rect 2134 2548 2138 2552
rect 2158 2548 2162 2552
rect 2054 2538 2058 2542
rect 2070 2538 2074 2542
rect 2038 2528 2042 2532
rect 2070 2528 2074 2532
rect 2030 2518 2034 2522
rect 2014 2498 2018 2502
rect 1990 2478 1994 2482
rect 2006 2478 2010 2482
rect 2038 2488 2042 2492
rect 1894 2458 1898 2462
rect 1958 2458 1962 2462
rect 1974 2458 1978 2462
rect 2006 2458 2010 2462
rect 1974 2448 1978 2452
rect 1982 2448 1986 2452
rect 2022 2448 2026 2452
rect 1910 2398 1914 2402
rect 2054 2468 2058 2472
rect 2102 2528 2106 2532
rect 2078 2508 2082 2512
rect 2094 2468 2098 2472
rect 2046 2458 2050 2462
rect 2070 2458 2074 2462
rect 2086 2448 2090 2452
rect 2038 2438 2042 2442
rect 2070 2438 2074 2442
rect 2030 2418 2034 2422
rect 1982 2388 1986 2392
rect 2006 2408 2010 2412
rect 2014 2408 2018 2412
rect 1910 2368 1914 2372
rect 1990 2368 1994 2372
rect 1854 2348 1858 2352
rect 2054 2368 2058 2372
rect 1950 2358 1954 2362
rect 1974 2358 1978 2362
rect 1942 2348 1946 2352
rect 2038 2348 2042 2352
rect 1854 2338 1858 2342
rect 1886 2338 1890 2342
rect 1966 2338 1970 2342
rect 1998 2338 2002 2342
rect 1870 2328 1874 2332
rect 1870 2308 1874 2312
rect 1878 2298 1882 2302
rect 1966 2328 1970 2332
rect 1966 2308 1970 2312
rect 1930 2303 1934 2307
rect 1937 2303 1941 2307
rect 1910 2298 1914 2302
rect 1838 2278 1842 2282
rect 1862 2278 1866 2282
rect 1902 2278 1906 2282
rect 1990 2298 1994 2302
rect 1974 2278 1978 2282
rect 1854 2258 1858 2262
rect 1814 2228 1818 2232
rect 1830 2228 1834 2232
rect 1758 2158 1762 2162
rect 1806 2158 1810 2162
rect 1830 2158 1834 2162
rect 1670 2148 1674 2152
rect 1718 2148 1722 2152
rect 1798 2148 1802 2152
rect 1870 2238 1874 2242
rect 1902 2258 1906 2262
rect 2022 2308 2026 2312
rect 2038 2308 2042 2312
rect 2030 2298 2034 2302
rect 2014 2268 2018 2272
rect 1918 2248 1922 2252
rect 1926 2248 1930 2252
rect 1942 2248 1946 2252
rect 1998 2258 2002 2262
rect 2030 2258 2034 2262
rect 1990 2248 1994 2252
rect 2014 2248 2018 2252
rect 2038 2248 2042 2252
rect 1918 2238 1922 2242
rect 1950 2238 1954 2242
rect 1910 2228 1914 2232
rect 1886 2208 1890 2212
rect 2078 2378 2082 2382
rect 2070 2338 2074 2342
rect 2062 2328 2066 2332
rect 1974 2228 1978 2232
rect 2046 2228 2050 2232
rect 2030 2218 2034 2222
rect 1966 2158 1970 2162
rect 1974 2158 1978 2162
rect 1910 2148 1914 2152
rect 2006 2148 2010 2152
rect 1646 2138 1650 2142
rect 1678 2138 1682 2142
rect 1702 2138 1706 2142
rect 1774 2138 1778 2142
rect 1846 2138 1850 2142
rect 1614 2118 1618 2122
rect 1614 2068 1618 2072
rect 1574 2058 1578 2062
rect 1590 2058 1594 2062
rect 1566 2048 1570 2052
rect 1550 1998 1554 2002
rect 1598 1998 1602 2002
rect 1646 2008 1650 2012
rect 1630 1988 1634 1992
rect 1574 1948 1578 1952
rect 1590 1938 1594 1942
rect 1566 1908 1570 1912
rect 1606 1908 1610 1912
rect 1686 2128 1690 2132
rect 1726 2128 1730 2132
rect 1758 2128 1762 2132
rect 1742 2118 1746 2122
rect 1806 2118 1810 2122
rect 1710 2098 1714 2102
rect 1758 2098 1762 2102
rect 1710 2088 1714 2092
rect 1726 2058 1730 2062
rect 1678 1988 1682 1992
rect 1734 1988 1738 1992
rect 1718 1968 1722 1972
rect 1718 1948 1722 1952
rect 1742 1948 1746 1952
rect 1678 1928 1682 1932
rect 1662 1918 1666 1922
rect 1670 1908 1674 1912
rect 1630 1898 1634 1902
rect 1662 1898 1666 1902
rect 1574 1888 1578 1892
rect 1614 1888 1618 1892
rect 1646 1888 1650 1892
rect 1494 1868 1498 1872
rect 1510 1868 1514 1872
rect 1534 1858 1538 1862
rect 1550 1858 1554 1862
rect 1566 1858 1570 1862
rect 1494 1838 1498 1842
rect 1550 1838 1554 1842
rect 1486 1808 1490 1812
rect 1582 1828 1586 1832
rect 1550 1778 1554 1782
rect 1430 1768 1434 1772
rect 1510 1768 1514 1772
rect 1534 1768 1538 1772
rect 1454 1758 1458 1762
rect 1518 1758 1522 1762
rect 1382 1748 1386 1752
rect 1414 1748 1418 1752
rect 1358 1738 1362 1742
rect 1326 1728 1330 1732
rect 1302 1688 1306 1692
rect 1310 1688 1314 1692
rect 1254 1678 1258 1682
rect 1278 1678 1282 1682
rect 1246 1668 1250 1672
rect 1214 1658 1218 1662
rect 1118 1648 1122 1652
rect 1038 1638 1042 1642
rect 1070 1638 1074 1642
rect 1094 1638 1098 1642
rect 1062 1608 1066 1612
rect 1070 1578 1074 1582
rect 1030 1558 1034 1562
rect 1070 1558 1074 1562
rect 1150 1628 1154 1632
rect 1102 1598 1106 1602
rect 1166 1598 1170 1602
rect 1198 1598 1202 1602
rect 1110 1588 1114 1592
rect 1134 1588 1138 1592
rect 1102 1578 1106 1582
rect 1182 1588 1186 1592
rect 1022 1548 1026 1552
rect 1014 1538 1018 1542
rect 1006 1518 1010 1522
rect 1014 1498 1018 1502
rect 1054 1548 1058 1552
rect 1086 1548 1090 1552
rect 1094 1548 1098 1552
rect 1054 1538 1058 1542
rect 1046 1518 1050 1522
rect 1046 1488 1050 1492
rect 1062 1488 1066 1492
rect 1070 1488 1074 1492
rect 1006 1458 1010 1462
rect 1086 1468 1090 1472
rect 1054 1458 1058 1462
rect 1038 1448 1042 1452
rect 1014 1438 1018 1442
rect 1022 1438 1026 1442
rect 1078 1418 1082 1422
rect 1006 1408 1010 1412
rect 1006 1368 1010 1372
rect 1046 1358 1050 1362
rect 1078 1358 1082 1362
rect 1118 1558 1122 1562
rect 1142 1558 1146 1562
rect 1190 1558 1194 1562
rect 1150 1548 1154 1552
rect 1126 1538 1130 1542
rect 1134 1518 1138 1522
rect 1198 1508 1202 1512
rect 1238 1658 1242 1662
rect 1238 1648 1242 1652
rect 1230 1638 1234 1642
rect 1262 1638 1266 1642
rect 1302 1628 1306 1632
rect 1278 1598 1282 1602
rect 1286 1598 1290 1602
rect 1222 1558 1226 1562
rect 1270 1558 1274 1562
rect 1278 1558 1282 1562
rect 1254 1548 1258 1552
rect 1342 1718 1346 1722
rect 1366 1718 1370 1722
rect 1398 1718 1402 1722
rect 1374 1708 1378 1712
rect 1390 1708 1394 1712
rect 1342 1688 1346 1692
rect 1318 1578 1322 1582
rect 1326 1578 1330 1582
rect 1302 1558 1306 1562
rect 1310 1558 1314 1562
rect 1294 1538 1298 1542
rect 1214 1528 1218 1532
rect 1262 1528 1266 1532
rect 1270 1528 1274 1532
rect 1206 1498 1210 1502
rect 1182 1488 1186 1492
rect 1222 1488 1226 1492
rect 1126 1448 1130 1452
rect 1118 1438 1122 1442
rect 1158 1418 1162 1422
rect 1150 1358 1154 1362
rect 1158 1358 1162 1362
rect 1054 1348 1058 1352
rect 1070 1348 1074 1352
rect 1094 1348 1098 1352
rect 1038 1338 1042 1342
rect 1118 1338 1122 1342
rect 1150 1338 1154 1342
rect 1022 1308 1026 1312
rect 998 1278 1002 1282
rect 982 1268 986 1272
rect 966 1218 970 1222
rect 806 1138 810 1142
rect 846 1138 850 1142
rect 902 1118 906 1122
rect 798 1078 802 1082
rect 862 1108 866 1112
rect 898 1103 902 1107
rect 905 1103 909 1107
rect 854 1088 858 1092
rect 902 1058 906 1062
rect 886 1008 890 1012
rect 782 988 786 992
rect 726 978 730 982
rect 702 938 706 942
rect 710 918 714 922
rect 678 908 682 912
rect 710 908 714 912
rect 678 878 682 882
rect 686 868 690 872
rect 654 858 658 862
rect 678 858 682 862
rect 718 878 722 882
rect 694 838 698 842
rect 686 818 690 822
rect 630 758 634 762
rect 646 728 650 732
rect 670 738 674 742
rect 662 728 666 732
rect 702 748 706 752
rect 934 1138 938 1142
rect 950 1148 954 1152
rect 950 1138 954 1142
rect 950 1118 954 1122
rect 942 1098 946 1102
rect 918 1028 922 1032
rect 950 1078 954 1082
rect 870 958 874 962
rect 894 958 898 962
rect 742 948 746 952
rect 806 948 810 952
rect 790 918 794 922
rect 790 908 794 912
rect 774 898 778 902
rect 758 878 762 882
rect 734 868 738 872
rect 798 878 802 882
rect 1022 1228 1026 1232
rect 990 1148 994 1152
rect 998 1148 1002 1152
rect 998 1138 1002 1142
rect 1022 1108 1026 1112
rect 1006 1088 1010 1092
rect 998 1078 1002 1082
rect 1014 1068 1018 1072
rect 902 938 906 942
rect 898 903 902 907
rect 905 903 909 907
rect 926 868 930 872
rect 758 858 762 862
rect 806 858 810 862
rect 830 858 834 862
rect 910 858 914 862
rect 758 848 762 852
rect 718 838 722 842
rect 726 818 730 822
rect 726 788 730 792
rect 718 768 722 772
rect 758 768 762 772
rect 774 758 778 762
rect 734 748 738 752
rect 750 748 754 752
rect 726 738 730 742
rect 710 728 714 732
rect 718 728 722 732
rect 654 708 658 712
rect 678 708 682 712
rect 590 698 594 702
rect 622 698 626 702
rect 630 688 634 692
rect 646 678 650 682
rect 622 588 626 592
rect 766 738 770 742
rect 766 678 770 682
rect 774 678 778 682
rect 718 668 722 672
rect 750 668 754 672
rect 710 648 714 652
rect 782 638 786 642
rect 630 578 634 582
rect 782 588 786 592
rect 990 1058 994 1062
rect 1006 1058 1010 1062
rect 1014 1008 1018 1012
rect 998 998 1002 1002
rect 974 948 978 952
rect 1054 1328 1058 1332
rect 1046 1268 1050 1272
rect 1038 1208 1042 1212
rect 1062 1178 1066 1182
rect 1030 1018 1034 1022
rect 1142 1328 1146 1332
rect 1086 1308 1090 1312
rect 1078 1288 1082 1292
rect 1182 1408 1186 1412
rect 1190 1398 1194 1402
rect 1206 1398 1210 1402
rect 1214 1398 1218 1402
rect 1182 1388 1186 1392
rect 1190 1378 1194 1382
rect 1198 1378 1202 1382
rect 1190 1348 1194 1352
rect 1166 1298 1170 1302
rect 1198 1288 1202 1292
rect 1102 1278 1106 1282
rect 1126 1278 1130 1282
rect 1182 1278 1186 1282
rect 1286 1518 1290 1522
rect 1294 1508 1298 1512
rect 1286 1448 1290 1452
rect 1270 1428 1274 1432
rect 1278 1428 1282 1432
rect 1270 1388 1274 1392
rect 1246 1358 1250 1362
rect 1230 1348 1234 1352
rect 1222 1338 1226 1342
rect 1262 1348 1266 1352
rect 1334 1528 1338 1532
rect 1358 1648 1362 1652
rect 1422 1698 1426 1702
rect 1414 1688 1418 1692
rect 1398 1678 1402 1682
rect 1382 1668 1386 1672
rect 1494 1748 1498 1752
rect 1590 1798 1594 1802
rect 1614 1778 1618 1782
rect 1646 1858 1650 1862
rect 1686 1878 1690 1882
rect 1638 1848 1642 1852
rect 1654 1848 1658 1852
rect 1670 1848 1674 1852
rect 1630 1828 1634 1832
rect 1630 1808 1634 1812
rect 1606 1748 1610 1752
rect 1622 1748 1626 1752
rect 1550 1738 1554 1742
rect 1526 1728 1530 1732
rect 1542 1728 1546 1732
rect 1558 1728 1562 1732
rect 1558 1718 1562 1722
rect 1494 1698 1498 1702
rect 1542 1698 1546 1702
rect 1446 1688 1450 1692
rect 1430 1678 1434 1682
rect 1494 1678 1498 1682
rect 1550 1678 1554 1682
rect 1454 1668 1458 1672
rect 1470 1668 1474 1672
rect 1534 1668 1538 1672
rect 1702 1908 1706 1912
rect 1742 1918 1746 1922
rect 1702 1868 1706 1872
rect 1726 1858 1730 1862
rect 1702 1848 1706 1852
rect 1694 1828 1698 1832
rect 1654 1798 1658 1802
rect 1758 1938 1762 1942
rect 1742 1858 1746 1862
rect 1734 1838 1738 1842
rect 1654 1778 1658 1782
rect 1838 2108 1842 2112
rect 1838 2088 1842 2092
rect 1846 2058 1850 2062
rect 1782 2038 1786 2042
rect 1822 2048 1826 2052
rect 1830 2008 1834 2012
rect 1846 2008 1850 2012
rect 1806 1988 1810 1992
rect 1838 1988 1842 1992
rect 1774 1968 1778 1972
rect 1798 1968 1802 1972
rect 1798 1948 1802 1952
rect 1782 1938 1786 1942
rect 1766 1918 1770 1922
rect 1774 1898 1778 1902
rect 1766 1888 1770 1892
rect 1758 1808 1762 1812
rect 1806 1928 1810 1932
rect 1798 1918 1802 1922
rect 1934 2138 1938 2142
rect 1950 2138 1954 2142
rect 1990 2138 1994 2142
rect 1998 2138 2002 2142
rect 1878 2078 1882 2082
rect 1870 2068 1874 2072
rect 1886 2068 1890 2072
rect 1930 2103 1934 2107
rect 1937 2103 1941 2107
rect 1950 2098 1954 2102
rect 1902 2068 1906 2072
rect 2150 2538 2154 2542
rect 2134 2508 2138 2512
rect 2126 2498 2130 2502
rect 2142 2498 2146 2502
rect 2134 2488 2138 2492
rect 2174 2528 2178 2532
rect 2158 2518 2162 2522
rect 2166 2518 2170 2522
rect 2174 2498 2178 2502
rect 2206 2648 2210 2652
rect 2198 2628 2202 2632
rect 2214 2598 2218 2602
rect 2246 2598 2250 2602
rect 2382 2658 2386 2662
rect 2414 2658 2418 2662
rect 2342 2648 2346 2652
rect 2366 2648 2370 2652
rect 2294 2638 2298 2642
rect 2326 2638 2330 2642
rect 2334 2628 2338 2632
rect 2278 2618 2282 2622
rect 2238 2588 2242 2592
rect 2326 2588 2330 2592
rect 2350 2598 2354 2602
rect 2342 2568 2346 2572
rect 2278 2558 2282 2562
rect 2230 2548 2234 2552
rect 2286 2548 2290 2552
rect 2198 2528 2202 2532
rect 2222 2528 2226 2532
rect 2222 2518 2226 2522
rect 2110 2428 2114 2432
rect 2126 2388 2130 2392
rect 2118 2368 2122 2372
rect 2142 2368 2146 2372
rect 2278 2538 2282 2542
rect 2318 2538 2322 2542
rect 2270 2528 2274 2532
rect 2254 2518 2258 2522
rect 2262 2508 2266 2512
rect 2246 2468 2250 2472
rect 2262 2468 2266 2472
rect 2214 2448 2218 2452
rect 2166 2428 2170 2432
rect 2158 2388 2162 2392
rect 2150 2358 2154 2362
rect 2302 2528 2306 2532
rect 2310 2528 2314 2532
rect 2294 2508 2298 2512
rect 2310 2498 2314 2502
rect 2302 2488 2306 2492
rect 2374 2628 2378 2632
rect 2422 2628 2426 2632
rect 2414 2608 2418 2612
rect 2398 2578 2402 2582
rect 2366 2548 2370 2552
rect 2510 2898 2514 2902
rect 2494 2828 2498 2832
rect 2502 2748 2506 2752
rect 2470 2668 2474 2672
rect 2462 2658 2466 2662
rect 2454 2638 2458 2642
rect 2442 2603 2446 2607
rect 2449 2603 2453 2607
rect 2422 2558 2426 2562
rect 2454 2558 2458 2562
rect 2334 2538 2338 2542
rect 2342 2528 2346 2532
rect 2430 2528 2434 2532
rect 2326 2458 2330 2462
rect 2294 2418 2298 2422
rect 2318 2418 2322 2422
rect 2278 2388 2282 2392
rect 2246 2378 2250 2382
rect 2206 2368 2210 2372
rect 2222 2368 2226 2372
rect 2174 2358 2178 2362
rect 2118 2348 2122 2352
rect 2166 2348 2170 2352
rect 2182 2348 2186 2352
rect 2206 2348 2210 2352
rect 2222 2348 2226 2352
rect 2238 2348 2242 2352
rect 2102 2338 2106 2342
rect 2094 2328 2098 2332
rect 2086 2318 2090 2322
rect 2094 2298 2098 2302
rect 2126 2338 2130 2342
rect 2214 2338 2218 2342
rect 2142 2308 2146 2312
rect 2078 2278 2082 2282
rect 2102 2278 2106 2282
rect 2142 2258 2146 2262
rect 2078 2248 2082 2252
rect 2094 2228 2098 2232
rect 2062 2198 2066 2202
rect 2070 2168 2074 2172
rect 2078 2168 2082 2172
rect 2038 2158 2042 2162
rect 2054 2158 2058 2162
rect 2046 2148 2050 2152
rect 2062 2148 2066 2152
rect 2046 2138 2050 2142
rect 2014 2128 2018 2132
rect 2054 2128 2058 2132
rect 1990 2098 1994 2102
rect 2022 2098 2026 2102
rect 1894 2058 1898 2062
rect 1974 2068 1978 2072
rect 1942 2048 1946 2052
rect 1870 2038 1874 2042
rect 1878 2038 1882 2042
rect 1862 2008 1866 2012
rect 1878 2008 1882 2012
rect 1894 2008 1898 2012
rect 1870 1988 1874 1992
rect 2038 2068 2042 2072
rect 2014 2048 2018 2052
rect 1998 2038 2002 2042
rect 2006 2038 2010 2042
rect 1966 1998 1970 2002
rect 1958 1988 1962 1992
rect 1926 1948 1930 1952
rect 1902 1938 1906 1942
rect 1974 1978 1978 1982
rect 1982 1968 1986 1972
rect 1998 1958 2002 1962
rect 2166 2168 2170 2172
rect 2110 2138 2114 2142
rect 2126 2138 2130 2142
rect 2094 2128 2098 2132
rect 2126 2118 2130 2122
rect 2062 2098 2066 2102
rect 2086 2088 2090 2092
rect 2078 2068 2082 2072
rect 2118 2068 2122 2072
rect 2126 2068 2130 2072
rect 2070 2058 2074 2062
rect 2110 2058 2114 2062
rect 2054 2048 2058 2052
rect 2038 2008 2042 2012
rect 2046 2008 2050 2012
rect 2014 1948 2018 1952
rect 1990 1938 1994 1942
rect 2014 1928 2018 1932
rect 2070 1998 2074 2002
rect 2038 1938 2042 1942
rect 1814 1908 1818 1912
rect 1854 1908 1858 1912
rect 1930 1903 1934 1907
rect 1937 1903 1941 1907
rect 1894 1898 1898 1902
rect 1870 1888 1874 1892
rect 1910 1888 1914 1892
rect 1918 1888 1922 1892
rect 1854 1848 1858 1852
rect 1790 1798 1794 1802
rect 1814 1798 1818 1802
rect 1734 1768 1738 1772
rect 1742 1768 1746 1772
rect 1774 1768 1778 1772
rect 1782 1768 1786 1772
rect 1678 1758 1682 1762
rect 1734 1758 1738 1762
rect 1670 1748 1674 1752
rect 1638 1738 1642 1742
rect 1598 1718 1602 1722
rect 1590 1708 1594 1712
rect 1654 1708 1658 1712
rect 1598 1698 1602 1702
rect 1646 1698 1650 1702
rect 1566 1688 1570 1692
rect 1574 1678 1578 1682
rect 1430 1658 1434 1662
rect 1462 1658 1466 1662
rect 1486 1658 1490 1662
rect 1502 1658 1506 1662
rect 1390 1648 1394 1652
rect 1374 1638 1378 1642
rect 1366 1598 1370 1602
rect 1358 1578 1362 1582
rect 1390 1598 1394 1602
rect 1418 1603 1422 1607
rect 1425 1603 1429 1607
rect 1454 1598 1458 1602
rect 1430 1558 1434 1562
rect 1358 1528 1362 1532
rect 1366 1518 1370 1522
rect 1342 1508 1346 1512
rect 1366 1508 1370 1512
rect 1390 1508 1394 1512
rect 1342 1498 1346 1502
rect 1350 1498 1354 1502
rect 1326 1488 1330 1492
rect 1310 1478 1314 1482
rect 1294 1358 1298 1362
rect 1398 1488 1402 1492
rect 1446 1528 1450 1532
rect 1438 1518 1442 1522
rect 1446 1508 1450 1512
rect 1358 1478 1362 1482
rect 1414 1478 1418 1482
rect 1342 1458 1346 1462
rect 1358 1458 1362 1462
rect 1318 1448 1322 1452
rect 1318 1398 1322 1402
rect 1390 1448 1394 1452
rect 1382 1438 1386 1442
rect 1374 1408 1378 1412
rect 1342 1388 1346 1392
rect 1342 1358 1346 1362
rect 1350 1358 1354 1362
rect 1446 1468 1450 1472
rect 1470 1598 1474 1602
rect 1502 1648 1506 1652
rect 1478 1568 1482 1572
rect 1486 1538 1490 1542
rect 1470 1498 1474 1502
rect 1622 1688 1626 1692
rect 1630 1678 1634 1682
rect 1726 1748 1730 1752
rect 1686 1738 1690 1742
rect 1710 1738 1714 1742
rect 1782 1748 1786 1752
rect 1694 1728 1698 1732
rect 1670 1688 1674 1692
rect 1662 1678 1666 1682
rect 1726 1688 1730 1692
rect 1750 1688 1754 1692
rect 1998 1918 2002 1922
rect 2030 1918 2034 1922
rect 1950 1868 1954 1872
rect 1958 1828 1962 1832
rect 1886 1728 1890 1732
rect 1782 1718 1786 1722
rect 1814 1718 1818 1722
rect 1870 1718 1874 1722
rect 1782 1678 1786 1682
rect 1710 1668 1714 1672
rect 1718 1668 1722 1672
rect 1614 1658 1618 1662
rect 1614 1648 1618 1652
rect 1590 1638 1594 1642
rect 1574 1608 1578 1612
rect 1566 1598 1570 1602
rect 1518 1588 1522 1592
rect 1510 1558 1514 1562
rect 1526 1568 1530 1572
rect 1566 1568 1570 1572
rect 1582 1568 1586 1572
rect 1542 1558 1546 1562
rect 1598 1628 1602 1632
rect 1622 1608 1626 1612
rect 1606 1568 1610 1572
rect 1614 1568 1618 1572
rect 1558 1548 1562 1552
rect 1646 1648 1650 1652
rect 1638 1608 1642 1612
rect 1550 1538 1554 1542
rect 1614 1538 1618 1542
rect 1630 1538 1634 1542
rect 1590 1528 1594 1532
rect 1470 1488 1474 1492
rect 1486 1488 1490 1492
rect 1526 1478 1530 1482
rect 1630 1528 1634 1532
rect 1638 1508 1642 1512
rect 1670 1638 1674 1642
rect 1710 1638 1714 1642
rect 1654 1538 1658 1542
rect 1718 1628 1722 1632
rect 1694 1608 1698 1612
rect 1678 1568 1682 1572
rect 1678 1558 1682 1562
rect 1670 1498 1674 1502
rect 1686 1498 1690 1502
rect 1686 1488 1690 1492
rect 1710 1508 1714 1512
rect 1710 1488 1714 1492
rect 1670 1478 1674 1482
rect 1702 1478 1706 1482
rect 1750 1648 1754 1652
rect 1774 1628 1778 1632
rect 1774 1608 1778 1612
rect 1774 1568 1778 1572
rect 1750 1558 1754 1562
rect 1758 1558 1762 1562
rect 1726 1548 1730 1552
rect 1750 1538 1754 1542
rect 1734 1498 1738 1502
rect 1766 1488 1770 1492
rect 1750 1478 1754 1482
rect 1502 1468 1506 1472
rect 1526 1468 1530 1472
rect 1574 1468 1578 1472
rect 1598 1468 1602 1472
rect 1686 1468 1690 1472
rect 1758 1468 1762 1472
rect 1446 1448 1450 1452
rect 1422 1438 1426 1442
rect 1438 1438 1442 1442
rect 1406 1408 1410 1412
rect 1418 1403 1422 1407
rect 1425 1403 1429 1407
rect 1390 1388 1394 1392
rect 1390 1378 1394 1382
rect 1414 1378 1418 1382
rect 1302 1348 1306 1352
rect 1318 1348 1322 1352
rect 1294 1338 1298 1342
rect 1230 1318 1234 1322
rect 1246 1318 1250 1322
rect 1230 1288 1234 1292
rect 1294 1318 1298 1322
rect 1286 1278 1290 1282
rect 1190 1268 1194 1272
rect 1270 1268 1274 1272
rect 1278 1268 1282 1272
rect 1094 1248 1098 1252
rect 1078 1238 1082 1242
rect 1326 1318 1330 1322
rect 1302 1268 1306 1272
rect 1310 1268 1314 1272
rect 1126 1258 1130 1262
rect 1158 1258 1162 1262
rect 1262 1258 1266 1262
rect 1182 1248 1186 1252
rect 1206 1248 1210 1252
rect 1102 1218 1106 1222
rect 1110 1178 1114 1182
rect 1070 1158 1074 1162
rect 1150 1238 1154 1242
rect 1166 1238 1170 1242
rect 1166 1218 1170 1222
rect 1246 1218 1250 1222
rect 1134 1208 1138 1212
rect 1158 1208 1162 1212
rect 1094 1158 1098 1162
rect 1118 1158 1122 1162
rect 1062 1148 1066 1152
rect 1078 1148 1082 1152
rect 1110 1148 1114 1152
rect 1126 1148 1130 1152
rect 1142 1158 1146 1162
rect 1086 1128 1090 1132
rect 1102 1128 1106 1132
rect 1054 1118 1058 1122
rect 1110 1108 1114 1112
rect 1070 1078 1074 1082
rect 1046 1058 1050 1062
rect 1054 1048 1058 1052
rect 1054 1028 1058 1032
rect 1078 1048 1082 1052
rect 1054 1008 1058 1012
rect 1070 1008 1074 1012
rect 1046 988 1050 992
rect 1022 978 1026 982
rect 1030 978 1034 982
rect 1038 978 1042 982
rect 1022 958 1026 962
rect 1006 948 1010 952
rect 1006 928 1010 932
rect 1022 918 1026 922
rect 982 878 986 882
rect 1014 878 1018 882
rect 1022 868 1026 872
rect 974 848 978 852
rect 966 838 970 842
rect 926 818 930 822
rect 870 808 874 812
rect 894 808 898 812
rect 838 728 842 732
rect 854 718 858 722
rect 878 708 882 712
rect 898 703 902 707
rect 905 703 909 707
rect 934 798 938 802
rect 934 778 938 782
rect 886 678 890 682
rect 814 668 818 672
rect 838 668 842 672
rect 1006 798 1010 802
rect 958 678 962 682
rect 822 658 826 662
rect 854 658 858 662
rect 950 658 954 662
rect 838 648 842 652
rect 806 588 810 592
rect 838 588 842 592
rect 798 568 802 572
rect 814 568 818 572
rect 926 648 930 652
rect 870 558 874 562
rect 582 548 586 552
rect 846 548 850 552
rect 862 548 866 552
rect 566 538 570 542
rect 486 408 490 412
rect 566 438 570 442
rect 558 428 562 432
rect 478 388 482 392
rect 526 388 530 392
rect 534 388 538 392
rect 390 268 394 272
rect 454 268 458 272
rect 414 258 418 262
rect 246 238 250 242
rect 358 228 362 232
rect 350 218 354 222
rect 318 188 322 192
rect 310 178 314 182
rect 214 148 218 152
rect 142 128 146 132
rect 230 118 234 122
rect 230 108 234 112
rect 166 98 170 102
rect 198 98 202 102
rect 30 78 34 82
rect 158 78 162 82
rect 342 158 346 162
rect 254 78 258 82
rect 6 48 10 52
rect 350 78 354 82
rect 342 68 346 72
rect 414 208 418 212
rect 394 203 398 207
rect 401 203 405 207
rect 374 68 378 72
rect 382 58 386 62
rect 326 28 330 32
rect 342 28 346 32
rect 358 8 362 12
rect 394 3 398 7
rect 401 3 405 7
rect 438 208 442 212
rect 574 398 578 402
rect 590 538 594 542
rect 526 348 530 352
rect 582 348 586 352
rect 710 528 714 532
rect 694 518 698 522
rect 694 498 698 502
rect 654 488 658 492
rect 806 538 810 542
rect 838 538 842 542
rect 758 518 762 522
rect 782 518 786 522
rect 750 498 754 502
rect 718 468 722 472
rect 742 468 746 472
rect 734 458 738 462
rect 670 438 674 442
rect 614 398 618 402
rect 686 388 690 392
rect 646 358 650 362
rect 678 358 682 362
rect 598 348 602 352
rect 614 348 618 352
rect 534 338 538 342
rect 590 338 594 342
rect 502 328 506 332
rect 582 298 586 302
rect 518 288 522 292
rect 534 288 538 292
rect 534 278 538 282
rect 630 298 634 302
rect 662 298 666 302
rect 694 338 698 342
rect 726 318 730 322
rect 670 278 674 282
rect 638 268 642 272
rect 614 228 618 232
rect 686 248 690 252
rect 614 218 618 222
rect 494 148 498 152
rect 582 148 586 152
rect 566 98 570 102
rect 526 88 530 92
rect 678 208 682 212
rect 630 148 634 152
rect 734 168 738 172
rect 694 148 698 152
rect 614 118 618 122
rect 438 58 442 62
rect 542 58 546 62
rect 582 58 586 62
rect 638 108 642 112
rect 638 78 642 82
rect 798 418 802 422
rect 782 398 786 402
rect 898 503 902 507
rect 905 503 909 507
rect 886 498 890 502
rect 862 488 866 492
rect 878 418 882 422
rect 822 398 826 402
rect 846 398 850 402
rect 814 378 818 382
rect 894 378 898 382
rect 934 608 938 612
rect 934 488 938 492
rect 814 348 818 352
rect 886 348 890 352
rect 902 348 906 352
rect 926 338 930 342
rect 854 328 858 332
rect 846 318 850 322
rect 758 298 762 302
rect 782 298 786 302
rect 774 288 778 292
rect 838 288 842 292
rect 898 303 902 307
rect 905 303 909 307
rect 806 278 810 282
rect 854 278 858 282
rect 814 268 818 272
rect 830 268 834 272
rect 790 198 794 202
rect 790 188 794 192
rect 766 98 770 102
rect 630 68 634 72
rect 678 58 682 62
rect 430 8 434 12
rect 446 8 450 12
rect 542 8 546 12
rect 558 8 562 12
rect 574 8 578 12
rect 630 8 634 12
rect 774 8 778 12
rect 822 258 826 262
rect 830 228 834 232
rect 830 178 834 182
rect 806 158 810 162
rect 822 158 826 162
rect 830 138 834 142
rect 918 268 922 272
rect 902 258 906 262
rect 862 248 866 252
rect 854 218 858 222
rect 878 208 882 212
rect 846 168 850 172
rect 894 228 898 232
rect 894 208 898 212
rect 902 208 906 212
rect 998 718 1002 722
rect 974 668 978 672
rect 1054 948 1058 952
rect 1070 948 1074 952
rect 1062 938 1066 942
rect 1038 848 1042 852
rect 1030 828 1034 832
rect 1070 928 1074 932
rect 1062 808 1066 812
rect 1094 998 1098 1002
rect 1094 938 1098 942
rect 1086 908 1090 912
rect 1110 958 1114 962
rect 1278 1138 1282 1142
rect 1310 1228 1314 1232
rect 1310 1198 1314 1202
rect 1302 1148 1306 1152
rect 1214 1128 1218 1132
rect 1294 1128 1298 1132
rect 1230 1118 1234 1122
rect 1166 1108 1170 1112
rect 1254 1108 1258 1112
rect 1278 1078 1282 1082
rect 1270 1068 1274 1072
rect 1326 1258 1330 1262
rect 1366 1338 1370 1342
rect 1422 1358 1426 1362
rect 1398 1338 1402 1342
rect 1422 1328 1426 1332
rect 1390 1298 1394 1302
rect 1342 1288 1346 1292
rect 1366 1288 1370 1292
rect 1366 1278 1370 1282
rect 1398 1278 1402 1282
rect 1342 1268 1346 1272
rect 1350 1268 1354 1272
rect 1374 1268 1378 1272
rect 1398 1258 1402 1262
rect 1358 1248 1362 1252
rect 1334 1188 1338 1192
rect 1342 1168 1346 1172
rect 1350 1168 1354 1172
rect 1326 1158 1330 1162
rect 1334 1158 1338 1162
rect 1318 1108 1322 1112
rect 1294 1058 1298 1062
rect 1278 1048 1282 1052
rect 1302 1048 1306 1052
rect 1174 1038 1178 1042
rect 1142 998 1146 1002
rect 1174 998 1178 1002
rect 1214 988 1218 992
rect 1198 958 1202 962
rect 1222 958 1226 962
rect 1126 948 1130 952
rect 1150 948 1154 952
rect 1182 948 1186 952
rect 1246 948 1250 952
rect 1262 948 1266 952
rect 1126 938 1130 942
rect 1142 938 1146 942
rect 1222 938 1226 942
rect 1238 938 1242 942
rect 1150 928 1154 932
rect 1166 918 1170 922
rect 1118 908 1122 912
rect 1134 888 1138 892
rect 1150 878 1154 882
rect 1262 928 1266 932
rect 1230 918 1234 922
rect 1262 918 1266 922
rect 1310 1038 1314 1042
rect 1286 948 1290 952
rect 1294 948 1298 952
rect 1294 928 1298 932
rect 1302 888 1306 892
rect 1286 878 1290 882
rect 1294 878 1298 882
rect 1102 808 1106 812
rect 1222 828 1226 832
rect 1206 778 1210 782
rect 1198 768 1202 772
rect 1126 758 1130 762
rect 1174 758 1178 762
rect 1214 758 1218 762
rect 1070 728 1074 732
rect 1078 728 1082 732
rect 1038 698 1042 702
rect 1118 738 1122 742
rect 1142 728 1146 732
rect 1174 738 1178 742
rect 1110 718 1114 722
rect 1150 718 1154 722
rect 1086 698 1090 702
rect 1134 698 1138 702
rect 1078 688 1082 692
rect 1110 678 1114 682
rect 1126 668 1130 672
rect 998 658 1002 662
rect 1022 658 1026 662
rect 1038 658 1042 662
rect 982 638 986 642
rect 1030 638 1034 642
rect 1014 618 1018 622
rect 966 598 970 602
rect 1086 588 1090 592
rect 998 578 1002 582
rect 982 568 986 572
rect 1086 558 1090 562
rect 1118 618 1122 622
rect 1046 548 1050 552
rect 1110 548 1114 552
rect 1214 738 1218 742
rect 1326 1078 1330 1082
rect 1334 1068 1338 1072
rect 1398 1248 1402 1252
rect 1446 1358 1450 1362
rect 1454 1348 1458 1352
rect 1462 1318 1466 1322
rect 1510 1458 1514 1462
rect 1510 1448 1514 1452
rect 1574 1458 1578 1462
rect 1582 1458 1586 1462
rect 1654 1458 1658 1462
rect 1750 1458 1754 1462
rect 1478 1378 1482 1382
rect 1502 1378 1506 1382
rect 1478 1348 1482 1352
rect 1486 1318 1490 1322
rect 1470 1308 1474 1312
rect 1462 1268 1466 1272
rect 1478 1268 1482 1272
rect 1494 1268 1498 1272
rect 1510 1268 1514 1272
rect 1454 1258 1458 1262
rect 1470 1258 1474 1262
rect 1422 1248 1426 1252
rect 1486 1248 1490 1252
rect 1406 1208 1410 1212
rect 1418 1203 1422 1207
rect 1425 1203 1429 1207
rect 1494 1198 1498 1202
rect 1438 1178 1442 1182
rect 1374 1158 1378 1162
rect 1422 1158 1426 1162
rect 1510 1228 1514 1232
rect 1558 1408 1562 1412
rect 1574 1408 1578 1412
rect 1558 1378 1562 1382
rect 1550 1358 1554 1362
rect 1526 1348 1530 1352
rect 1550 1338 1554 1342
rect 1542 1308 1546 1312
rect 1526 1298 1530 1302
rect 1534 1298 1538 1302
rect 1534 1278 1538 1282
rect 1526 1268 1530 1272
rect 1542 1248 1546 1252
rect 1550 1248 1554 1252
rect 1654 1448 1658 1452
rect 1590 1398 1594 1402
rect 1638 1398 1642 1402
rect 1654 1398 1658 1402
rect 1606 1388 1610 1392
rect 1622 1358 1626 1362
rect 1646 1358 1650 1362
rect 1574 1338 1578 1342
rect 1566 1318 1570 1322
rect 1574 1308 1578 1312
rect 1614 1318 1618 1322
rect 1566 1268 1570 1272
rect 1566 1238 1570 1242
rect 1566 1198 1570 1202
rect 1510 1188 1514 1192
rect 1574 1178 1578 1182
rect 1446 1148 1450 1152
rect 1462 1148 1466 1152
rect 1350 1108 1354 1112
rect 1358 1108 1362 1112
rect 1350 1088 1354 1092
rect 1374 1118 1378 1122
rect 1366 1078 1370 1082
rect 1382 1108 1386 1112
rect 1422 1108 1426 1112
rect 1406 1088 1410 1092
rect 1430 1098 1434 1102
rect 1382 1058 1386 1062
rect 1462 1138 1466 1142
rect 1486 1138 1490 1142
rect 1502 1128 1506 1132
rect 1478 1118 1482 1122
rect 1502 1118 1506 1122
rect 1510 1118 1514 1122
rect 1462 1098 1466 1102
rect 1446 1088 1450 1092
rect 1438 1068 1442 1072
rect 1406 1058 1410 1062
rect 1350 1048 1354 1052
rect 1390 1048 1394 1052
rect 1390 1008 1394 1012
rect 1374 998 1378 1002
rect 1342 978 1346 982
rect 1326 968 1330 972
rect 1358 958 1362 962
rect 1418 1003 1422 1007
rect 1425 1003 1429 1007
rect 1478 1068 1482 1072
rect 1526 1128 1530 1132
rect 1542 1128 1546 1132
rect 1630 1348 1634 1352
rect 1638 1318 1642 1322
rect 1670 1388 1674 1392
rect 1654 1268 1658 1272
rect 1622 1258 1626 1262
rect 1614 1248 1618 1252
rect 1606 1208 1610 1212
rect 1622 1218 1626 1222
rect 1598 1168 1602 1172
rect 1582 1158 1586 1162
rect 1566 1128 1570 1132
rect 1582 1118 1586 1122
rect 1590 1118 1594 1122
rect 1606 1118 1610 1122
rect 1518 1098 1522 1102
rect 1550 1098 1554 1102
rect 1510 1088 1514 1092
rect 1534 1088 1538 1092
rect 1550 1088 1554 1092
rect 1574 1088 1578 1092
rect 1574 1078 1578 1082
rect 1526 1068 1530 1072
rect 1534 1068 1538 1072
rect 1550 1068 1554 1072
rect 1478 1058 1482 1062
rect 1510 1058 1514 1062
rect 1614 1098 1618 1102
rect 1638 1198 1642 1202
rect 1702 1438 1706 1442
rect 1686 1428 1690 1432
rect 1726 1388 1730 1392
rect 1718 1378 1722 1382
rect 1694 1348 1698 1352
rect 1702 1318 1706 1322
rect 1686 1298 1690 1302
rect 1670 1258 1674 1262
rect 1678 1238 1682 1242
rect 1670 1198 1674 1202
rect 1662 1188 1666 1192
rect 1654 1168 1658 1172
rect 1630 1128 1634 1132
rect 1646 1118 1650 1122
rect 1638 1088 1642 1092
rect 1622 1078 1626 1082
rect 1646 1078 1650 1082
rect 1582 1058 1586 1062
rect 1606 1048 1610 1052
rect 1542 1038 1546 1042
rect 1470 1018 1474 1022
rect 1534 1008 1538 1012
rect 1446 958 1450 962
rect 1478 958 1482 962
rect 1502 958 1506 962
rect 1534 958 1538 962
rect 1350 948 1354 952
rect 1374 948 1378 952
rect 1342 928 1346 932
rect 1318 898 1322 902
rect 1326 898 1330 902
rect 1326 888 1330 892
rect 1342 888 1346 892
rect 1310 878 1314 882
rect 1350 878 1354 882
rect 1430 938 1434 942
rect 1382 928 1386 932
rect 1366 918 1370 922
rect 1406 888 1410 892
rect 1486 948 1490 952
rect 1478 938 1482 942
rect 1486 938 1490 942
rect 1510 938 1514 942
rect 1478 928 1482 932
rect 1462 918 1466 922
rect 1454 908 1458 912
rect 1454 888 1458 892
rect 1358 868 1362 872
rect 1310 858 1314 862
rect 1310 838 1314 842
rect 1270 818 1274 822
rect 1286 808 1290 812
rect 1366 858 1370 862
rect 1366 848 1370 852
rect 1374 838 1378 842
rect 1390 848 1394 852
rect 1350 798 1354 802
rect 1326 788 1330 792
rect 1262 778 1266 782
rect 1254 758 1258 762
rect 1462 868 1466 872
rect 1462 858 1466 862
rect 1478 858 1482 862
rect 1430 818 1434 822
rect 1418 803 1422 807
rect 1425 803 1429 807
rect 1406 798 1410 802
rect 1422 788 1426 792
rect 1470 768 1474 772
rect 1526 928 1530 932
rect 1494 908 1498 912
rect 1526 898 1530 902
rect 1502 888 1506 892
rect 1494 838 1498 842
rect 1486 808 1490 812
rect 1478 758 1482 762
rect 1510 868 1514 872
rect 1510 838 1514 842
rect 1494 758 1498 762
rect 1302 748 1306 752
rect 1462 748 1466 752
rect 1350 738 1354 742
rect 1470 738 1474 742
rect 1486 738 1490 742
rect 1246 728 1250 732
rect 1318 728 1322 732
rect 1238 708 1242 712
rect 1198 698 1202 702
rect 1238 698 1242 702
rect 1294 698 1298 702
rect 1246 688 1250 692
rect 1238 668 1242 672
rect 1278 668 1282 672
rect 1166 658 1170 662
rect 1214 658 1218 662
rect 1214 648 1218 652
rect 1230 648 1234 652
rect 1246 648 1250 652
rect 1262 648 1266 652
rect 1334 688 1338 692
rect 1286 658 1290 662
rect 1310 658 1314 662
rect 1462 728 1466 732
rect 1494 728 1498 732
rect 1390 708 1394 712
rect 1374 678 1378 682
rect 1382 678 1386 682
rect 1310 648 1314 652
rect 1270 628 1274 632
rect 1198 618 1202 622
rect 1334 618 1338 622
rect 1142 598 1146 602
rect 1126 558 1130 562
rect 1158 548 1162 552
rect 1278 548 1282 552
rect 1126 528 1130 532
rect 982 518 986 522
rect 974 508 978 512
rect 1070 498 1074 502
rect 1014 488 1018 492
rect 1046 488 1050 492
rect 990 478 994 482
rect 982 468 986 472
rect 982 458 986 462
rect 950 398 954 402
rect 942 358 946 362
rect 974 368 978 372
rect 966 348 970 352
rect 1022 448 1026 452
rect 1078 488 1082 492
rect 1118 488 1122 492
rect 1230 538 1234 542
rect 1166 518 1170 522
rect 1142 488 1146 492
rect 1134 478 1138 482
rect 1310 578 1314 582
rect 1326 558 1330 562
rect 1430 708 1434 712
rect 1398 698 1402 702
rect 1446 688 1450 692
rect 1438 678 1442 682
rect 1454 678 1458 682
rect 1430 668 1434 672
rect 1446 668 1450 672
rect 1494 708 1498 712
rect 1502 708 1506 712
rect 1470 678 1474 682
rect 1486 678 1490 682
rect 1494 678 1498 682
rect 1478 668 1482 672
rect 1494 668 1498 672
rect 1454 658 1458 662
rect 1358 578 1362 582
rect 1374 578 1378 582
rect 1382 578 1386 582
rect 1302 518 1306 522
rect 1270 488 1274 492
rect 1214 478 1218 482
rect 1254 478 1258 482
rect 1110 468 1114 472
rect 1142 468 1146 472
rect 1182 468 1186 472
rect 990 438 994 442
rect 1054 438 1058 442
rect 1014 418 1018 422
rect 998 378 1002 382
rect 1062 408 1066 412
rect 1102 438 1106 442
rect 1030 398 1034 402
rect 1094 398 1098 402
rect 1046 358 1050 362
rect 1070 358 1074 362
rect 1094 358 1098 362
rect 982 318 986 322
rect 1030 348 1034 352
rect 1054 338 1058 342
rect 1062 338 1066 342
rect 1086 338 1090 342
rect 1086 318 1090 322
rect 1014 298 1018 302
rect 1046 268 1050 272
rect 1166 458 1170 462
rect 1126 448 1130 452
rect 1142 448 1146 452
rect 1134 388 1138 392
rect 1142 368 1146 372
rect 1190 368 1194 372
rect 1190 358 1194 362
rect 1150 348 1154 352
rect 1182 348 1186 352
rect 1198 348 1202 352
rect 1094 298 1098 302
rect 950 258 954 262
rect 1030 258 1034 262
rect 934 188 938 192
rect 966 248 970 252
rect 1030 218 1034 222
rect 950 208 954 212
rect 942 178 946 182
rect 966 168 970 172
rect 1014 168 1018 172
rect 894 158 898 162
rect 934 158 938 162
rect 942 158 946 162
rect 982 158 986 162
rect 846 148 850 152
rect 902 148 906 152
rect 982 148 986 152
rect 1014 148 1018 152
rect 1062 198 1066 202
rect 1038 168 1042 172
rect 1054 168 1058 172
rect 958 138 962 142
rect 990 138 994 142
rect 1022 138 1026 142
rect 1038 138 1042 142
rect 1126 338 1130 342
rect 1150 328 1154 332
rect 1118 278 1122 282
rect 1134 278 1138 282
rect 1310 448 1314 452
rect 1222 408 1226 412
rect 1294 408 1298 412
rect 1238 368 1242 372
rect 1286 368 1290 372
rect 1262 358 1266 362
rect 1230 338 1234 342
rect 1214 318 1218 322
rect 1238 318 1242 322
rect 1198 298 1202 302
rect 1422 638 1426 642
rect 1422 618 1426 622
rect 1390 568 1394 572
rect 1418 603 1422 607
rect 1425 603 1429 607
rect 1438 598 1442 602
rect 1390 548 1394 552
rect 1406 548 1410 552
rect 1414 548 1418 552
rect 1446 568 1450 572
rect 1462 648 1466 652
rect 1494 648 1498 652
rect 1486 638 1490 642
rect 1454 548 1458 552
rect 1478 548 1482 552
rect 1430 538 1434 542
rect 1374 528 1378 532
rect 1398 528 1402 532
rect 1414 478 1418 482
rect 1358 468 1362 472
rect 1382 458 1386 462
rect 1334 448 1338 452
rect 1326 378 1330 382
rect 1318 368 1322 372
rect 1390 438 1394 442
rect 1358 418 1362 422
rect 1350 368 1354 372
rect 1358 368 1362 372
rect 1374 368 1378 372
rect 1318 358 1322 362
rect 1334 358 1338 362
rect 1350 338 1354 342
rect 1286 328 1290 332
rect 1310 328 1314 332
rect 1270 298 1274 302
rect 1334 298 1338 302
rect 1174 278 1178 282
rect 1230 278 1234 282
rect 1318 278 1322 282
rect 1182 268 1186 272
rect 1214 268 1218 272
rect 1278 268 1282 272
rect 1294 268 1298 272
rect 1118 258 1122 262
rect 1110 218 1114 222
rect 1094 208 1098 212
rect 1078 188 1082 192
rect 1086 188 1090 192
rect 1198 258 1202 262
rect 1206 258 1210 262
rect 1214 248 1218 252
rect 1166 238 1170 242
rect 1158 228 1162 232
rect 1086 168 1090 172
rect 1110 168 1114 172
rect 1078 158 1082 162
rect 1230 228 1234 232
rect 1166 188 1170 192
rect 1190 188 1194 192
rect 1214 188 1218 192
rect 1134 158 1138 162
rect 1126 138 1130 142
rect 1142 138 1146 142
rect 1150 138 1154 142
rect 814 108 818 112
rect 838 88 842 92
rect 806 68 810 72
rect 806 58 810 62
rect 862 128 866 132
rect 998 128 1002 132
rect 1070 128 1074 132
rect 1086 128 1090 132
rect 1118 128 1122 132
rect 1134 128 1138 132
rect 878 118 882 122
rect 870 108 874 112
rect 1038 108 1042 112
rect 854 88 858 92
rect 898 103 902 107
rect 905 103 909 107
rect 942 88 946 92
rect 918 78 922 82
rect 870 68 874 72
rect 910 68 914 72
rect 870 58 874 62
rect 934 58 938 62
rect 998 78 1002 82
rect 1030 78 1034 82
rect 974 68 978 72
rect 1022 68 1026 72
rect 1118 78 1122 82
rect 1086 68 1090 72
rect 1110 68 1114 72
rect 1014 58 1018 62
rect 1038 58 1042 62
rect 878 48 882 52
rect 1030 48 1034 52
rect 1062 48 1066 52
rect 1190 168 1194 172
rect 1262 228 1266 232
rect 1254 188 1258 192
rect 1238 178 1242 182
rect 1246 178 1250 182
rect 1238 168 1242 172
rect 1230 158 1234 162
rect 1262 158 1266 162
rect 1198 138 1202 142
rect 1246 138 1250 142
rect 1174 88 1178 92
rect 1230 88 1234 92
rect 1174 68 1178 72
rect 1302 258 1306 262
rect 1294 248 1298 252
rect 1310 248 1314 252
rect 1382 338 1386 342
rect 1374 268 1378 272
rect 1382 268 1386 272
rect 1350 248 1354 252
rect 1350 228 1354 232
rect 1358 228 1362 232
rect 1310 218 1314 222
rect 1318 188 1322 192
rect 1302 158 1306 162
rect 1334 178 1338 182
rect 1326 158 1330 162
rect 1334 158 1338 162
rect 1310 138 1314 142
rect 1286 128 1290 132
rect 1318 128 1322 132
rect 1366 208 1370 212
rect 1478 528 1482 532
rect 1462 498 1466 502
rect 1454 478 1458 482
rect 1590 1028 1594 1032
rect 1598 1028 1602 1032
rect 1574 1008 1578 1012
rect 1670 1158 1674 1162
rect 1670 1118 1674 1122
rect 1710 1308 1714 1312
rect 1710 1268 1714 1272
rect 1742 1348 1746 1352
rect 1734 1318 1738 1322
rect 1750 1318 1754 1322
rect 1734 1308 1738 1312
rect 1702 1258 1706 1262
rect 1694 1148 1698 1152
rect 1694 1118 1698 1122
rect 1930 1703 1934 1707
rect 1937 1703 1941 1707
rect 1830 1698 1834 1702
rect 1862 1698 1866 1702
rect 1854 1688 1858 1692
rect 1918 1688 1922 1692
rect 1934 1688 1938 1692
rect 1822 1678 1826 1682
rect 1838 1678 1842 1682
rect 1870 1678 1874 1682
rect 1790 1648 1794 1652
rect 1798 1638 1802 1642
rect 1814 1638 1818 1642
rect 1886 1648 1890 1652
rect 1862 1628 1866 1632
rect 1854 1618 1858 1622
rect 1814 1608 1818 1612
rect 1838 1568 1842 1572
rect 1790 1558 1794 1562
rect 1798 1548 1802 1552
rect 1806 1548 1810 1552
rect 1830 1548 1834 1552
rect 1838 1548 1842 1552
rect 1918 1648 1922 1652
rect 1926 1648 1930 1652
rect 1910 1618 1914 1622
rect 1942 1638 1946 1642
rect 1934 1608 1938 1612
rect 2054 1908 2058 1912
rect 2022 1898 2026 1902
rect 2006 1878 2010 1882
rect 2054 1878 2058 1882
rect 2022 1868 2026 1872
rect 1990 1818 1994 1822
rect 1958 1768 1962 1772
rect 1982 1768 1986 1772
rect 2030 1858 2034 1862
rect 2054 1858 2058 1862
rect 2094 1878 2098 1882
rect 2094 1858 2098 1862
rect 2086 1848 2090 1852
rect 2078 1818 2082 1822
rect 2070 1808 2074 1812
rect 2078 1798 2082 1802
rect 2230 2328 2234 2332
rect 2254 2318 2258 2322
rect 2262 2298 2266 2302
rect 2230 2248 2234 2252
rect 2182 2198 2186 2202
rect 2174 2128 2178 2132
rect 2158 2108 2162 2112
rect 2150 2098 2154 2102
rect 2214 2188 2218 2192
rect 2214 2168 2218 2172
rect 2214 2158 2218 2162
rect 2198 2148 2202 2152
rect 2158 2058 2162 2062
rect 2126 2048 2130 2052
rect 2142 2048 2146 2052
rect 2230 2108 2234 2112
rect 2262 2138 2266 2142
rect 2302 2368 2306 2372
rect 2350 2518 2354 2522
rect 2366 2518 2370 2522
rect 2382 2498 2386 2502
rect 2374 2458 2378 2462
rect 2486 2638 2490 2642
rect 2502 2608 2506 2612
rect 2510 2598 2514 2602
rect 2486 2588 2490 2592
rect 2486 2568 2490 2572
rect 2462 2518 2466 2522
rect 2398 2478 2402 2482
rect 2390 2448 2394 2452
rect 2406 2448 2410 2452
rect 2358 2438 2362 2442
rect 2350 2408 2354 2412
rect 2414 2438 2418 2442
rect 2494 2558 2498 2562
rect 2542 2988 2546 2992
rect 2526 2878 2530 2882
rect 2954 3103 2958 3107
rect 2961 3103 2965 3107
rect 3978 3103 3982 3107
rect 3985 3103 3989 3107
rect 2638 3098 2642 3102
rect 3614 3088 3618 3092
rect 3646 3088 3650 3092
rect 3862 3088 3866 3092
rect 4094 3088 4098 3092
rect 4262 3088 4266 3092
rect 3054 3078 3058 3082
rect 3502 3078 3506 3082
rect 3558 3078 3562 3082
rect 3590 3078 3594 3082
rect 2670 3068 2674 3072
rect 2606 3058 2610 3062
rect 2662 3058 2666 3062
rect 2606 3028 2610 3032
rect 2726 3058 2730 3062
rect 2670 3008 2674 3012
rect 2566 2978 2570 2982
rect 2566 2968 2570 2972
rect 2750 2998 2754 3002
rect 2814 2998 2818 3002
rect 2766 2968 2770 2972
rect 2798 2968 2802 2972
rect 2726 2958 2730 2962
rect 2598 2948 2602 2952
rect 2654 2948 2658 2952
rect 2758 2948 2762 2952
rect 2558 2928 2562 2932
rect 2798 2928 2802 2932
rect 2806 2928 2810 2932
rect 2566 2918 2570 2922
rect 2582 2918 2586 2922
rect 2670 2918 2674 2922
rect 2742 2918 2746 2922
rect 2782 2918 2786 2922
rect 2902 3058 2906 3062
rect 2950 3058 2954 3062
rect 2870 2968 2874 2972
rect 2862 2958 2866 2962
rect 2838 2928 2842 2932
rect 2822 2898 2826 2902
rect 2830 2898 2834 2902
rect 2846 2918 2850 2922
rect 2550 2878 2554 2882
rect 2574 2878 2578 2882
rect 2614 2878 2618 2882
rect 2630 2878 2634 2882
rect 2814 2878 2818 2882
rect 2526 2858 2530 2862
rect 2534 2848 2538 2852
rect 2566 2768 2570 2772
rect 2542 2748 2546 2752
rect 2534 2738 2538 2742
rect 2526 2698 2530 2702
rect 2502 2548 2506 2552
rect 2478 2508 2482 2512
rect 2510 2498 2514 2502
rect 2598 2858 2602 2862
rect 2590 2818 2594 2822
rect 2590 2768 2594 2772
rect 2638 2848 2642 2852
rect 2606 2818 2610 2822
rect 2670 2808 2674 2812
rect 2870 2948 2874 2952
rect 2886 2918 2890 2922
rect 2998 3018 3002 3022
rect 2902 2978 2906 2982
rect 2974 2958 2978 2962
rect 2910 2948 2914 2952
rect 2998 2948 3002 2952
rect 2910 2928 2914 2932
rect 2942 2918 2946 2922
rect 2902 2898 2906 2902
rect 2894 2878 2898 2882
rect 2838 2868 2842 2872
rect 2862 2858 2866 2862
rect 2750 2788 2754 2792
rect 2622 2768 2626 2772
rect 2662 2768 2666 2772
rect 2750 2768 2754 2772
rect 2582 2748 2586 2752
rect 2598 2748 2602 2752
rect 2574 2738 2578 2742
rect 2566 2728 2570 2732
rect 2598 2718 2602 2722
rect 2542 2708 2546 2712
rect 2582 2708 2586 2712
rect 2542 2698 2546 2702
rect 2622 2698 2626 2702
rect 2534 2678 2538 2682
rect 2582 2688 2586 2692
rect 2598 2688 2602 2692
rect 2582 2668 2586 2672
rect 2558 2568 2562 2572
rect 2662 2748 2666 2752
rect 2694 2748 2698 2752
rect 2654 2738 2658 2742
rect 2686 2738 2690 2742
rect 2718 2738 2722 2742
rect 2726 2728 2730 2732
rect 2702 2708 2706 2712
rect 2694 2698 2698 2702
rect 2678 2678 2682 2682
rect 2734 2678 2738 2682
rect 2798 2748 2802 2752
rect 2830 2748 2834 2752
rect 2750 2738 2754 2742
rect 2782 2738 2786 2742
rect 2806 2738 2810 2742
rect 2758 2728 2762 2732
rect 2774 2728 2778 2732
rect 2750 2718 2754 2722
rect 2790 2718 2794 2722
rect 2846 2728 2850 2732
rect 2838 2708 2842 2712
rect 2830 2698 2834 2702
rect 2710 2668 2714 2672
rect 2718 2668 2722 2672
rect 2742 2668 2746 2672
rect 2750 2668 2754 2672
rect 2638 2658 2642 2662
rect 2638 2648 2642 2652
rect 2670 2648 2674 2652
rect 2686 2648 2690 2652
rect 2670 2638 2674 2642
rect 2590 2558 2594 2562
rect 2654 2548 2658 2552
rect 2534 2538 2538 2542
rect 2550 2538 2554 2542
rect 2542 2518 2546 2522
rect 2574 2518 2578 2522
rect 2606 2538 2610 2542
rect 2622 2528 2626 2532
rect 2654 2528 2658 2532
rect 2766 2658 2770 2662
rect 2742 2648 2746 2652
rect 2750 2648 2754 2652
rect 2702 2638 2706 2642
rect 2718 2618 2722 2622
rect 2718 2598 2722 2602
rect 2798 2648 2802 2652
rect 2814 2618 2818 2622
rect 2790 2578 2794 2582
rect 2718 2558 2722 2562
rect 2670 2518 2674 2522
rect 2614 2508 2618 2512
rect 2662 2508 2666 2512
rect 2702 2518 2706 2522
rect 2598 2498 2602 2502
rect 2502 2488 2506 2492
rect 2486 2468 2490 2472
rect 2574 2478 2578 2482
rect 2606 2478 2610 2482
rect 2630 2488 2634 2492
rect 2630 2478 2634 2482
rect 2582 2468 2586 2472
rect 2606 2468 2610 2472
rect 2590 2458 2594 2462
rect 2646 2458 2650 2462
rect 2446 2448 2450 2452
rect 2486 2448 2490 2452
rect 2614 2448 2618 2452
rect 2442 2403 2446 2407
rect 2449 2403 2453 2407
rect 2430 2398 2434 2402
rect 2502 2438 2506 2442
rect 2414 2378 2418 2382
rect 2342 2348 2346 2352
rect 2358 2348 2362 2352
rect 2342 2338 2346 2342
rect 2390 2338 2394 2342
rect 2342 2318 2346 2322
rect 2366 2298 2370 2302
rect 2334 2268 2338 2272
rect 2350 2268 2354 2272
rect 2398 2278 2402 2282
rect 2566 2418 2570 2422
rect 2542 2368 2546 2372
rect 2566 2368 2570 2372
rect 2478 2358 2482 2362
rect 2518 2358 2522 2362
rect 2462 2348 2466 2352
rect 2478 2348 2482 2352
rect 2710 2498 2714 2502
rect 2694 2488 2698 2492
rect 2774 2548 2778 2552
rect 2790 2528 2794 2532
rect 2774 2498 2778 2502
rect 2734 2478 2738 2482
rect 2886 2748 2890 2752
rect 2878 2738 2882 2742
rect 2862 2698 2866 2702
rect 2954 2903 2958 2907
rect 2961 2903 2965 2907
rect 2950 2858 2954 2862
rect 2982 2858 2986 2862
rect 2934 2828 2938 2832
rect 3006 2818 3010 2822
rect 3086 3058 3090 3062
rect 3118 3058 3122 3062
rect 3054 3038 3058 3042
rect 3102 3028 3106 3032
rect 3118 2948 3122 2952
rect 3070 2938 3074 2942
rect 3102 2918 3106 2922
rect 3054 2898 3058 2902
rect 3078 2898 3082 2902
rect 3110 2898 3114 2902
rect 3126 2888 3130 2892
rect 3094 2878 3098 2882
rect 3230 3058 3234 3062
rect 3294 3058 3298 3062
rect 3190 3038 3194 3042
rect 3198 3018 3202 3022
rect 3206 2968 3210 2972
rect 3142 2948 3146 2952
rect 3158 2948 3162 2952
rect 3166 2938 3170 2942
rect 3142 2848 3146 2852
rect 2998 2798 3002 2802
rect 3014 2798 3018 2802
rect 3062 2798 3066 2802
rect 3134 2798 3138 2802
rect 2918 2788 2922 2792
rect 2918 2768 2922 2772
rect 3014 2768 3018 2772
rect 3102 2768 3106 2772
rect 3190 2948 3194 2952
rect 3270 2988 3274 2992
rect 3294 2958 3298 2962
rect 3222 2948 3226 2952
rect 3206 2928 3210 2932
rect 3190 2898 3194 2902
rect 3198 2858 3202 2862
rect 3278 2928 3282 2932
rect 3278 2918 3282 2922
rect 3366 3048 3370 3052
rect 3518 3058 3522 3062
rect 3566 3058 3570 3062
rect 3678 3078 3682 3082
rect 3750 3078 3754 3082
rect 3766 3078 3770 3082
rect 3854 3078 3858 3082
rect 3886 3078 3890 3082
rect 4150 3078 4154 3082
rect 4182 3078 4186 3082
rect 4286 3078 4290 3082
rect 3694 3068 3698 3072
rect 3622 3058 3626 3062
rect 3550 3048 3554 3052
rect 3614 3048 3618 3052
rect 3494 3038 3498 3042
rect 3526 3038 3530 3042
rect 3454 3018 3458 3022
rect 3474 3003 3478 3007
rect 3481 3003 3485 3007
rect 3558 3028 3562 3032
rect 3566 3028 3570 3032
rect 3502 3008 3506 3012
rect 3518 3008 3522 3012
rect 3558 2988 3562 2992
rect 3422 2958 3426 2962
rect 3438 2958 3442 2962
rect 3446 2958 3450 2962
rect 3478 2958 3482 2962
rect 3494 2958 3498 2962
rect 3406 2948 3410 2952
rect 3430 2948 3434 2952
rect 3478 2948 3482 2952
rect 3438 2938 3442 2942
rect 3382 2928 3386 2932
rect 3414 2928 3418 2932
rect 3366 2918 3370 2922
rect 3374 2908 3378 2912
rect 3318 2898 3322 2902
rect 3334 2898 3338 2902
rect 3350 2898 3354 2902
rect 3230 2878 3234 2882
rect 3278 2878 3282 2882
rect 3246 2858 3250 2862
rect 3270 2858 3274 2862
rect 3350 2858 3354 2862
rect 3190 2848 3194 2852
rect 3214 2848 3218 2852
rect 3262 2848 3266 2852
rect 3254 2828 3258 2832
rect 3174 2798 3178 2802
rect 3566 2978 3570 2982
rect 3502 2918 3506 2922
rect 3550 2908 3554 2912
rect 3502 2898 3506 2902
rect 3534 2898 3538 2902
rect 3478 2888 3482 2892
rect 3494 2888 3498 2892
rect 3518 2888 3522 2892
rect 3526 2888 3530 2892
rect 3502 2878 3506 2882
rect 3454 2818 3458 2822
rect 3406 2808 3410 2812
rect 3446 2808 3450 2812
rect 3366 2788 3370 2792
rect 3166 2778 3170 2782
rect 3326 2778 3330 2782
rect 3430 2768 3434 2772
rect 3446 2768 3450 2772
rect 3542 2878 3546 2882
rect 3558 2878 3562 2882
rect 3670 3058 3674 3062
rect 3702 3058 3706 3062
rect 3686 3048 3690 3052
rect 3742 3068 3746 3072
rect 3790 3068 3794 3072
rect 3822 3068 3826 3072
rect 3758 3058 3762 3062
rect 3766 3048 3770 3052
rect 3782 3048 3786 3052
rect 3798 3048 3802 3052
rect 3654 3038 3658 3042
rect 3670 3038 3674 3042
rect 3702 3038 3706 3042
rect 3718 3038 3722 3042
rect 3670 3028 3674 3032
rect 3606 3018 3610 3022
rect 3654 3018 3658 3022
rect 3582 2978 3586 2982
rect 3718 3008 3722 3012
rect 3710 2998 3714 3002
rect 3670 2988 3674 2992
rect 3614 2958 3618 2962
rect 3622 2958 3626 2962
rect 3638 2958 3642 2962
rect 3694 2978 3698 2982
rect 3654 2948 3658 2952
rect 3718 2988 3722 2992
rect 3766 3038 3770 3042
rect 3774 3038 3778 3042
rect 3766 2978 3770 2982
rect 3742 2968 3746 2972
rect 3758 2968 3762 2972
rect 3830 3048 3834 3052
rect 3822 3038 3826 3042
rect 3814 3008 3818 3012
rect 3822 2988 3826 2992
rect 3830 2988 3834 2992
rect 3798 2968 3802 2972
rect 3782 2958 3786 2962
rect 3590 2928 3594 2932
rect 3678 2928 3682 2932
rect 3686 2928 3690 2932
rect 3702 2928 3706 2932
rect 3734 2928 3738 2932
rect 3574 2888 3578 2892
rect 3638 2918 3642 2922
rect 3630 2898 3634 2902
rect 3598 2878 3602 2882
rect 3494 2858 3498 2862
rect 3550 2858 3554 2862
rect 3574 2858 3578 2862
rect 3494 2848 3498 2852
rect 3518 2848 3522 2852
rect 3494 2808 3498 2812
rect 3474 2803 3478 2807
rect 3481 2803 3485 2807
rect 3510 2788 3514 2792
rect 3470 2768 3474 2772
rect 3542 2838 3546 2842
rect 3550 2798 3554 2802
rect 3574 2838 3578 2842
rect 3566 2788 3570 2792
rect 3598 2858 3602 2862
rect 3614 2858 3618 2862
rect 3590 2818 3594 2822
rect 3566 2758 3570 2762
rect 3582 2758 3586 2762
rect 3086 2748 3090 2752
rect 3126 2748 3130 2752
rect 3134 2748 3138 2752
rect 3166 2748 3170 2752
rect 3222 2748 3226 2752
rect 3382 2748 3386 2752
rect 3398 2748 3402 2752
rect 3446 2748 3450 2752
rect 3518 2748 3522 2752
rect 2958 2728 2962 2732
rect 2910 2718 2914 2722
rect 2998 2718 3002 2722
rect 2954 2703 2958 2707
rect 2961 2703 2965 2707
rect 3046 2698 3050 2702
rect 3014 2678 3018 2682
rect 3030 2678 3034 2682
rect 2838 2618 2842 2622
rect 2854 2608 2858 2612
rect 2846 2548 2850 2552
rect 2814 2488 2818 2492
rect 2678 2468 2682 2472
rect 2694 2468 2698 2472
rect 2742 2468 2746 2472
rect 2798 2468 2802 2472
rect 2814 2468 2818 2472
rect 2686 2428 2690 2432
rect 2734 2458 2738 2462
rect 2750 2458 2754 2462
rect 2758 2448 2762 2452
rect 2750 2428 2754 2432
rect 2766 2428 2770 2432
rect 2678 2388 2682 2392
rect 2654 2378 2658 2382
rect 2582 2368 2586 2372
rect 2606 2368 2610 2372
rect 2630 2368 2634 2372
rect 2654 2368 2658 2372
rect 2662 2368 2666 2372
rect 2782 2448 2786 2452
rect 2790 2408 2794 2412
rect 2774 2388 2778 2392
rect 2766 2368 2770 2372
rect 2806 2378 2810 2382
rect 2774 2358 2778 2362
rect 2798 2358 2802 2362
rect 2590 2348 2594 2352
rect 2742 2348 2746 2352
rect 2854 2448 2858 2452
rect 2846 2418 2850 2422
rect 2838 2398 2842 2402
rect 2822 2388 2826 2392
rect 2950 2668 2954 2672
rect 2998 2668 3002 2672
rect 3030 2668 3034 2672
rect 3062 2668 3066 2672
rect 3110 2738 3114 2742
rect 3134 2738 3138 2742
rect 3094 2728 3098 2732
rect 3118 2708 3122 2712
rect 3238 2738 3242 2742
rect 3086 2688 3090 2692
rect 3102 2688 3106 2692
rect 3094 2668 3098 2672
rect 3110 2668 3114 2672
rect 3022 2658 3026 2662
rect 3070 2658 3074 2662
rect 3118 2658 3122 2662
rect 3254 2708 3258 2712
rect 3262 2688 3266 2692
rect 3406 2738 3410 2742
rect 3358 2718 3362 2722
rect 3414 2728 3418 2732
rect 3494 2728 3498 2732
rect 3398 2718 3402 2722
rect 3462 2718 3466 2722
rect 3382 2708 3386 2712
rect 3502 2708 3506 2712
rect 3286 2688 3290 2692
rect 3430 2688 3434 2692
rect 3166 2678 3170 2682
rect 3190 2678 3194 2682
rect 3278 2678 3282 2682
rect 3366 2678 3370 2682
rect 3166 2668 3170 2672
rect 3278 2668 3282 2672
rect 3310 2668 3314 2672
rect 3166 2658 3170 2662
rect 3134 2648 3138 2652
rect 3150 2648 3154 2652
rect 3062 2638 3066 2642
rect 3086 2638 3090 2642
rect 3110 2638 3114 2642
rect 2918 2608 2922 2612
rect 3054 2578 3058 2582
rect 3030 2558 3034 2562
rect 2910 2548 2914 2552
rect 2966 2548 2970 2552
rect 3006 2538 3010 2542
rect 2910 2528 2914 2532
rect 2902 2508 2906 2512
rect 2950 2518 2954 2522
rect 2934 2508 2938 2512
rect 2926 2478 2930 2482
rect 2870 2458 2874 2462
rect 2910 2458 2914 2462
rect 2894 2438 2898 2442
rect 2870 2378 2874 2382
rect 2918 2448 2922 2452
rect 2954 2503 2958 2507
rect 2961 2503 2965 2507
rect 2958 2488 2962 2492
rect 2982 2468 2986 2472
rect 3006 2468 3010 2472
rect 3174 2638 3178 2642
rect 3142 2628 3146 2632
rect 3110 2608 3114 2612
rect 3086 2578 3090 2582
rect 3150 2568 3154 2572
rect 3150 2548 3154 2552
rect 3038 2458 3042 2462
rect 2950 2418 2954 2422
rect 2998 2418 3002 2422
rect 2974 2398 2978 2402
rect 3030 2408 3034 2412
rect 3022 2378 3026 2382
rect 2910 2368 2914 2372
rect 3014 2368 3018 2372
rect 2862 2358 2866 2362
rect 2878 2358 2882 2362
rect 2902 2358 2906 2362
rect 2814 2348 2818 2352
rect 2846 2348 2850 2352
rect 2878 2348 2882 2352
rect 2454 2338 2458 2342
rect 2518 2338 2522 2342
rect 2526 2338 2530 2342
rect 2574 2338 2578 2342
rect 2638 2338 2642 2342
rect 2678 2338 2682 2342
rect 2750 2338 2754 2342
rect 2790 2338 2794 2342
rect 2446 2318 2450 2322
rect 2470 2308 2474 2312
rect 2454 2278 2458 2282
rect 2390 2268 2394 2272
rect 2422 2268 2426 2272
rect 2446 2268 2450 2272
rect 2318 2258 2322 2262
rect 2342 2258 2346 2262
rect 2382 2238 2386 2242
rect 2302 2198 2306 2202
rect 2278 2188 2282 2192
rect 2366 2188 2370 2192
rect 2326 2178 2330 2182
rect 2318 2168 2322 2172
rect 2366 2158 2370 2162
rect 2294 2148 2298 2152
rect 2286 2138 2290 2142
rect 2334 2138 2338 2142
rect 2350 2138 2354 2142
rect 2270 2128 2274 2132
rect 2334 2128 2338 2132
rect 2286 2098 2290 2102
rect 2318 2098 2322 2102
rect 2246 2088 2250 2092
rect 2390 2198 2394 2202
rect 2442 2203 2446 2207
rect 2449 2203 2453 2207
rect 2534 2328 2538 2332
rect 2566 2328 2570 2332
rect 2574 2318 2578 2322
rect 2550 2308 2554 2312
rect 2494 2278 2498 2282
rect 2558 2268 2562 2272
rect 2510 2248 2514 2252
rect 2486 2238 2490 2242
rect 2502 2198 2506 2202
rect 2478 2178 2482 2182
rect 2414 2158 2418 2162
rect 2446 2148 2450 2152
rect 2486 2148 2490 2152
rect 2382 2128 2386 2132
rect 2358 2108 2362 2112
rect 2430 2128 2434 2132
rect 2406 2108 2410 2112
rect 2382 2098 2386 2102
rect 2398 2098 2402 2102
rect 2614 2298 2618 2302
rect 2582 2268 2586 2272
rect 2606 2268 2610 2272
rect 2574 2258 2578 2262
rect 2590 2258 2594 2262
rect 2566 2228 2570 2232
rect 2574 2228 2578 2232
rect 2526 2178 2530 2182
rect 2550 2178 2554 2182
rect 2534 2138 2538 2142
rect 2438 2108 2442 2112
rect 2382 2078 2386 2082
rect 2414 2078 2418 2082
rect 2462 2128 2466 2132
rect 2542 2128 2546 2132
rect 2470 2098 2474 2102
rect 2502 2078 2506 2082
rect 2526 2098 2530 2102
rect 2694 2328 2698 2332
rect 2710 2328 2714 2332
rect 2766 2328 2770 2332
rect 2838 2338 2842 2342
rect 2926 2358 2930 2362
rect 3006 2358 3010 2362
rect 2886 2338 2890 2342
rect 2894 2338 2898 2342
rect 2854 2328 2858 2332
rect 2822 2318 2826 2322
rect 2830 2318 2834 2322
rect 2750 2308 2754 2312
rect 2998 2348 3002 2352
rect 2934 2338 2938 2342
rect 2990 2338 2994 2342
rect 3022 2338 3026 2342
rect 2974 2328 2978 2332
rect 2954 2303 2958 2307
rect 2961 2303 2965 2307
rect 2662 2278 2666 2282
rect 2942 2278 2946 2282
rect 2734 2268 2738 2272
rect 2638 2248 2642 2252
rect 2638 2218 2642 2222
rect 2646 2218 2650 2222
rect 2622 2208 2626 2212
rect 2566 2148 2570 2152
rect 2574 2138 2578 2142
rect 2590 2138 2594 2142
rect 2558 2118 2562 2122
rect 2694 2198 2698 2202
rect 2654 2148 2658 2152
rect 2678 2148 2682 2152
rect 2718 2188 2722 2192
rect 2726 2178 2730 2182
rect 2734 2148 2738 2152
rect 2654 2138 2658 2142
rect 2686 2138 2690 2142
rect 2630 2128 2634 2132
rect 2686 2118 2690 2122
rect 2598 2108 2602 2112
rect 2638 2098 2642 2102
rect 2646 2098 2650 2102
rect 2622 2088 2626 2092
rect 2550 2078 2554 2082
rect 2422 2068 2426 2072
rect 2438 2068 2442 2072
rect 2510 2068 2514 2072
rect 2302 2058 2306 2062
rect 2350 2058 2354 2062
rect 2366 2058 2370 2062
rect 2206 2008 2210 2012
rect 2198 1998 2202 2002
rect 2414 2058 2418 2062
rect 2494 2058 2498 2062
rect 2510 2058 2514 2062
rect 2478 2028 2482 2032
rect 2398 2008 2402 2012
rect 2442 2003 2446 2007
rect 2449 2003 2453 2007
rect 2534 2048 2538 2052
rect 2550 2048 2554 2052
rect 2582 2048 2586 2052
rect 2534 2028 2538 2032
rect 2478 1958 2482 1962
rect 2510 1958 2514 1962
rect 2166 1948 2170 1952
rect 2278 1948 2282 1952
rect 2366 1948 2370 1952
rect 2382 1948 2386 1952
rect 2486 1948 2490 1952
rect 2502 1948 2506 1952
rect 2518 1948 2522 1952
rect 2166 1938 2170 1942
rect 2230 1938 2234 1942
rect 2326 1938 2330 1942
rect 2366 1938 2370 1942
rect 2222 1928 2226 1932
rect 2246 1928 2250 1932
rect 2182 1918 2186 1922
rect 2134 1908 2138 1912
rect 2126 1898 2130 1902
rect 2118 1888 2122 1892
rect 2182 1888 2186 1892
rect 2278 1918 2282 1922
rect 2262 1908 2266 1912
rect 2214 1878 2218 1882
rect 2230 1878 2234 1882
rect 2198 1868 2202 1872
rect 2142 1858 2146 1862
rect 2166 1848 2170 1852
rect 2262 1866 2266 1870
rect 2246 1858 2250 1862
rect 2174 1798 2178 1802
rect 2062 1778 2066 1782
rect 2110 1778 2114 1782
rect 2182 1778 2186 1782
rect 2070 1768 2074 1772
rect 2054 1758 2058 1762
rect 2078 1758 2082 1762
rect 1982 1738 1986 1742
rect 1998 1738 2002 1742
rect 1990 1728 1994 1732
rect 1958 1698 1962 1702
rect 1958 1618 1962 1622
rect 2158 1768 2162 1772
rect 2150 1758 2154 1762
rect 2190 1758 2194 1762
rect 2062 1748 2066 1752
rect 2070 1738 2074 1742
rect 2022 1728 2026 1732
rect 2030 1728 2034 1732
rect 2046 1728 2050 1732
rect 2006 1708 2010 1712
rect 2022 1708 2026 1712
rect 1998 1698 2002 1702
rect 2014 1698 2018 1702
rect 2022 1678 2026 1682
rect 2038 1708 2042 1712
rect 2054 1698 2058 1702
rect 2222 1848 2226 1852
rect 2254 1848 2258 1852
rect 2454 1918 2458 1922
rect 2462 1918 2466 1922
rect 2294 1908 2298 1912
rect 2358 1908 2362 1912
rect 2414 1908 2418 1912
rect 2430 1908 2434 1912
rect 2302 1888 2306 1892
rect 2294 1858 2298 1862
rect 2382 1888 2386 1892
rect 2398 1888 2402 1892
rect 2334 1868 2338 1872
rect 2318 1858 2322 1862
rect 2278 1808 2282 1812
rect 2222 1758 2226 1762
rect 2238 1758 2242 1762
rect 2270 1758 2274 1762
rect 2342 1848 2346 1852
rect 2326 1818 2330 1822
rect 2366 1858 2370 1862
rect 2382 1858 2386 1862
rect 2406 1868 2410 1872
rect 2406 1838 2410 1842
rect 2390 1818 2394 1822
rect 2358 1768 2362 1772
rect 2438 1898 2442 1902
rect 2430 1878 2434 1882
rect 2502 1908 2506 1912
rect 2534 1928 2538 1932
rect 2510 1868 2514 1872
rect 2478 1858 2482 1862
rect 2502 1858 2506 1862
rect 2574 2028 2578 2032
rect 2558 1968 2562 1972
rect 2614 2008 2618 2012
rect 2646 2008 2650 2012
rect 2662 1988 2666 1992
rect 2582 1978 2586 1982
rect 2622 1968 2626 1972
rect 2590 1958 2594 1962
rect 2630 1958 2634 1962
rect 2598 1938 2602 1942
rect 2662 1938 2666 1942
rect 2566 1918 2570 1922
rect 2686 1928 2690 1932
rect 2654 1898 2658 1902
rect 2590 1888 2594 1892
rect 2678 1888 2682 1892
rect 2606 1878 2610 1882
rect 2678 1868 2682 1872
rect 2542 1858 2546 1862
rect 2662 1858 2666 1862
rect 2534 1838 2538 1842
rect 2502 1818 2506 1822
rect 2526 1818 2530 1822
rect 2442 1803 2446 1807
rect 2449 1803 2453 1807
rect 2478 1768 2482 1772
rect 2486 1768 2490 1772
rect 2310 1748 2314 1752
rect 2462 1748 2466 1752
rect 2158 1738 2162 1742
rect 2182 1738 2186 1742
rect 2198 1738 2202 1742
rect 2214 1738 2218 1742
rect 2086 1728 2090 1732
rect 2102 1728 2106 1732
rect 2118 1728 2122 1732
rect 2110 1688 2114 1692
rect 2134 1708 2138 1712
rect 2246 1738 2250 1742
rect 2230 1728 2234 1732
rect 2270 1718 2274 1722
rect 2142 1698 2146 1702
rect 2126 1678 2130 1682
rect 2278 1708 2282 1712
rect 2246 1698 2250 1702
rect 2262 1688 2266 1692
rect 2126 1668 2130 1672
rect 2150 1668 2154 1672
rect 2022 1658 2026 1662
rect 2062 1658 2066 1662
rect 2086 1658 2090 1662
rect 2110 1658 2114 1662
rect 1998 1648 2002 1652
rect 2070 1648 2074 1652
rect 1974 1628 1978 1632
rect 1998 1628 2002 1632
rect 2062 1618 2066 1622
rect 2094 1608 2098 1612
rect 1950 1588 1954 1592
rect 1862 1558 1866 1562
rect 1950 1558 1954 1562
rect 1870 1548 1874 1552
rect 1902 1548 1906 1552
rect 1894 1538 1898 1542
rect 1846 1508 1850 1512
rect 1942 1538 1946 1542
rect 1894 1518 1898 1522
rect 1822 1478 1826 1482
rect 1838 1478 1842 1482
rect 1814 1468 1818 1472
rect 1830 1468 1834 1472
rect 1782 1458 1786 1462
rect 1822 1458 1826 1462
rect 1854 1458 1858 1462
rect 1798 1448 1802 1452
rect 1830 1448 1834 1452
rect 1774 1388 1778 1392
rect 1766 1358 1770 1362
rect 1766 1348 1770 1352
rect 1814 1348 1818 1352
rect 1782 1318 1786 1322
rect 1806 1318 1810 1322
rect 1854 1398 1858 1402
rect 1846 1388 1850 1392
rect 1870 1448 1874 1452
rect 1878 1388 1882 1392
rect 1886 1358 1890 1362
rect 2086 1598 2090 1602
rect 2006 1588 2010 1592
rect 2022 1588 2026 1592
rect 2054 1588 2058 1592
rect 1982 1558 1986 1562
rect 1966 1548 1970 1552
rect 1998 1548 2002 1552
rect 1958 1518 1962 1522
rect 1930 1503 1934 1507
rect 1937 1503 1941 1507
rect 2030 1558 2034 1562
rect 2022 1538 2026 1542
rect 1974 1488 1978 1492
rect 1926 1478 1930 1482
rect 2046 1518 2050 1522
rect 2174 1668 2178 1672
rect 2358 1738 2362 1742
rect 2374 1728 2378 1732
rect 2478 1708 2482 1712
rect 2382 1688 2386 1692
rect 2142 1638 2146 1642
rect 2166 1638 2170 1642
rect 2278 1638 2282 1642
rect 2118 1568 2122 1572
rect 2158 1558 2162 1562
rect 2118 1548 2122 1552
rect 2158 1548 2162 1552
rect 2094 1538 2098 1542
rect 2102 1540 2106 1542
rect 2102 1538 2106 1540
rect 2118 1538 2122 1542
rect 2070 1508 2074 1512
rect 2038 1498 2042 1502
rect 1902 1468 1906 1472
rect 2070 1468 2074 1472
rect 1910 1458 1914 1462
rect 1974 1458 1978 1462
rect 1998 1458 2002 1462
rect 2014 1458 2018 1462
rect 1918 1398 1922 1402
rect 1902 1378 1906 1382
rect 1846 1348 1850 1352
rect 1854 1348 1858 1352
rect 1870 1348 1874 1352
rect 1894 1348 1898 1352
rect 1902 1338 1906 1342
rect 1838 1328 1842 1332
rect 1854 1318 1858 1322
rect 1886 1318 1890 1322
rect 1830 1308 1834 1312
rect 1790 1298 1794 1302
rect 1814 1298 1818 1302
rect 1814 1288 1818 1292
rect 1766 1268 1770 1272
rect 1742 1188 1746 1192
rect 1734 1168 1738 1172
rect 1718 1138 1722 1142
rect 1750 1168 1754 1172
rect 1766 1218 1770 1222
rect 1822 1268 1826 1272
rect 1782 1258 1786 1262
rect 1798 1258 1802 1262
rect 1830 1258 1834 1262
rect 1886 1308 1890 1312
rect 1878 1278 1882 1282
rect 1774 1198 1778 1202
rect 1854 1228 1858 1232
rect 1814 1188 1818 1192
rect 1894 1298 1898 1302
rect 1902 1268 1906 1272
rect 1910 1248 1914 1252
rect 1910 1218 1914 1222
rect 2022 1448 2026 1452
rect 1990 1438 1994 1442
rect 1974 1418 1978 1422
rect 1958 1368 1962 1372
rect 1958 1358 1962 1362
rect 1958 1348 1962 1352
rect 1926 1328 1930 1332
rect 1950 1328 1954 1332
rect 1930 1303 1934 1307
rect 1937 1303 1941 1307
rect 1958 1268 1962 1272
rect 1942 1258 1946 1262
rect 1918 1188 1922 1192
rect 1878 1178 1882 1182
rect 1942 1178 1946 1182
rect 1838 1168 1842 1172
rect 1790 1148 1794 1152
rect 1822 1148 1826 1152
rect 1718 1128 1722 1132
rect 1750 1128 1754 1132
rect 1822 1128 1826 1132
rect 1830 1128 1834 1132
rect 1702 1098 1706 1102
rect 1734 1098 1738 1102
rect 1686 1078 1690 1082
rect 1662 1058 1666 1062
rect 1646 1048 1650 1052
rect 1638 1038 1642 1042
rect 1574 978 1578 982
rect 1638 958 1642 962
rect 1582 948 1586 952
rect 1550 908 1554 912
rect 1542 888 1546 892
rect 1542 878 1546 882
rect 1558 898 1562 902
rect 1542 868 1546 872
rect 1598 938 1602 942
rect 1582 908 1586 912
rect 1582 888 1586 892
rect 1574 868 1578 872
rect 1638 928 1642 932
rect 1614 918 1618 922
rect 1614 898 1618 902
rect 1582 838 1586 842
rect 1686 1048 1690 1052
rect 1710 1078 1714 1082
rect 1774 1088 1778 1092
rect 1694 998 1698 1002
rect 1694 988 1698 992
rect 1670 958 1674 962
rect 1718 978 1722 982
rect 1726 958 1730 962
rect 1702 948 1706 952
rect 1646 878 1650 882
rect 1638 868 1642 872
rect 1598 828 1602 832
rect 1638 798 1642 802
rect 1590 788 1594 792
rect 1622 778 1626 782
rect 1558 768 1562 772
rect 1574 768 1578 772
rect 1598 768 1602 772
rect 1526 758 1530 762
rect 1542 758 1546 762
rect 1526 728 1530 732
rect 1518 718 1522 722
rect 1526 718 1530 722
rect 1630 748 1634 752
rect 1574 718 1578 722
rect 1566 698 1570 702
rect 1566 678 1570 682
rect 1518 658 1522 662
rect 1502 628 1506 632
rect 1526 638 1530 642
rect 1518 628 1522 632
rect 1638 738 1642 742
rect 1622 728 1626 732
rect 1630 728 1634 732
rect 1606 708 1610 712
rect 1742 938 1746 942
rect 1662 858 1666 862
rect 1662 838 1666 842
rect 1670 828 1674 832
rect 1702 888 1706 892
rect 1742 918 1746 922
rect 1718 898 1722 902
rect 1726 888 1730 892
rect 1734 878 1738 882
rect 1686 868 1690 872
rect 1710 868 1714 872
rect 1694 858 1698 862
rect 1702 858 1706 862
rect 1726 858 1730 862
rect 1678 808 1682 812
rect 1686 768 1690 772
rect 1702 838 1706 842
rect 1734 808 1738 812
rect 1702 798 1706 802
rect 1726 758 1730 762
rect 1726 748 1730 752
rect 1670 738 1674 742
rect 1686 738 1690 742
rect 1702 738 1706 742
rect 1662 718 1666 722
rect 1638 708 1642 712
rect 1646 708 1650 712
rect 1654 708 1658 712
rect 1654 698 1658 702
rect 1726 718 1730 722
rect 1702 678 1706 682
rect 1606 668 1610 672
rect 1614 658 1618 662
rect 1678 658 1682 662
rect 1590 638 1594 642
rect 1590 608 1594 612
rect 1502 568 1506 572
rect 1510 568 1514 572
rect 1534 568 1538 572
rect 1614 558 1618 562
rect 1670 648 1674 652
rect 1654 638 1658 642
rect 1638 618 1642 622
rect 1630 568 1634 572
rect 1646 608 1650 612
rect 1502 548 1506 552
rect 1534 548 1538 552
rect 1566 548 1570 552
rect 1598 548 1602 552
rect 1518 528 1522 532
rect 1550 528 1554 532
rect 1510 508 1514 512
rect 1550 498 1554 502
rect 1478 478 1482 482
rect 1510 478 1514 482
rect 1534 478 1538 482
rect 1478 468 1482 472
rect 1494 468 1498 472
rect 1454 458 1458 462
rect 1462 458 1466 462
rect 1478 458 1482 462
rect 1418 403 1422 407
rect 1425 403 1429 407
rect 1398 378 1402 382
rect 1486 398 1490 402
rect 1454 368 1458 372
rect 1422 358 1426 362
rect 1470 358 1474 362
rect 1398 268 1402 272
rect 1438 268 1442 272
rect 1382 258 1386 262
rect 1406 258 1410 262
rect 1430 258 1434 262
rect 1438 228 1442 232
rect 1382 218 1386 222
rect 1422 218 1426 222
rect 1418 203 1422 207
rect 1425 203 1429 207
rect 1398 198 1402 202
rect 1390 158 1394 162
rect 1374 138 1378 142
rect 1326 108 1330 112
rect 1366 128 1370 132
rect 1382 118 1386 122
rect 1358 98 1362 102
rect 1526 468 1530 472
rect 1534 448 1538 452
rect 1510 368 1514 372
rect 1510 358 1514 362
rect 1526 358 1530 362
rect 1470 338 1474 342
rect 1494 338 1498 342
rect 1526 338 1530 342
rect 1518 328 1522 332
rect 1462 318 1466 322
rect 1486 318 1490 322
rect 1494 308 1498 312
rect 1518 278 1522 282
rect 1542 338 1546 342
rect 1542 328 1546 332
rect 1534 278 1538 282
rect 1502 268 1506 272
rect 1526 268 1530 272
rect 1590 538 1594 542
rect 1606 528 1610 532
rect 1598 518 1602 522
rect 1590 478 1594 482
rect 1566 468 1570 472
rect 1582 468 1586 472
rect 1606 468 1610 472
rect 1646 538 1650 542
rect 1622 528 1626 532
rect 1662 568 1666 572
rect 1814 1078 1818 1082
rect 1822 1078 1826 1082
rect 1854 1158 1858 1162
rect 1878 1158 1882 1162
rect 1894 1158 1898 1162
rect 1846 1138 1850 1142
rect 1878 1138 1882 1142
rect 1862 1128 1866 1132
rect 1846 1098 1850 1102
rect 1878 1098 1882 1102
rect 1870 1088 1874 1092
rect 1862 1078 1866 1082
rect 1790 1068 1794 1072
rect 1806 1068 1810 1072
rect 1982 1388 1986 1392
rect 1990 1338 1994 1342
rect 2062 1448 2066 1452
rect 2038 1398 2042 1402
rect 2038 1388 2042 1392
rect 2046 1378 2050 1382
rect 2006 1358 2010 1362
rect 2022 1358 2026 1362
rect 2054 1358 2058 1362
rect 2062 1358 2066 1362
rect 2054 1338 2058 1342
rect 2094 1448 2098 1452
rect 2094 1418 2098 1422
rect 1998 1328 2002 1332
rect 2030 1308 2034 1312
rect 2078 1308 2082 1312
rect 1990 1278 1994 1282
rect 2070 1298 2074 1302
rect 2222 1618 2226 1622
rect 2214 1608 2218 1612
rect 2198 1568 2202 1572
rect 2286 1598 2290 1602
rect 2270 1568 2274 1572
rect 2182 1548 2186 1552
rect 2134 1528 2138 1532
rect 2174 1528 2178 1532
rect 2182 1528 2186 1532
rect 2134 1518 2138 1522
rect 2294 1558 2298 1562
rect 2246 1548 2250 1552
rect 2262 1538 2266 1542
rect 2262 1518 2266 1522
rect 2230 1488 2234 1492
rect 2230 1478 2234 1482
rect 2118 1468 2122 1472
rect 2214 1468 2218 1472
rect 2110 1458 2114 1462
rect 2302 1458 2306 1462
rect 2214 1438 2218 1442
rect 2126 1428 2130 1432
rect 2110 1378 2114 1382
rect 2102 1358 2106 1362
rect 2310 1448 2314 1452
rect 2366 1658 2370 1662
rect 2358 1558 2362 1562
rect 2374 1538 2378 1542
rect 2350 1518 2354 1522
rect 2334 1498 2338 1502
rect 2326 1468 2330 1472
rect 2334 1458 2338 1462
rect 2374 1458 2378 1462
rect 2358 1448 2362 1452
rect 2310 1428 2314 1432
rect 2286 1378 2290 1382
rect 2342 1388 2346 1392
rect 2358 1388 2362 1392
rect 2318 1378 2322 1382
rect 2302 1358 2306 1362
rect 2286 1348 2290 1352
rect 2302 1348 2306 1352
rect 2326 1358 2330 1362
rect 2342 1348 2346 1352
rect 2534 1758 2538 1762
rect 2502 1688 2506 1692
rect 2398 1678 2402 1682
rect 2398 1658 2402 1662
rect 2710 2118 2714 2122
rect 2806 2258 2810 2262
rect 2854 2258 2858 2262
rect 2886 2258 2890 2262
rect 2822 2218 2826 2222
rect 2838 2218 2842 2222
rect 2926 2248 2930 2252
rect 2910 2188 2914 2192
rect 2894 2178 2898 2182
rect 2822 2148 2826 2152
rect 3046 2378 3050 2382
rect 3062 2508 3066 2512
rect 3102 2518 3106 2522
rect 3142 2538 3146 2542
rect 3158 2538 3162 2542
rect 3166 2538 3170 2542
rect 3126 2498 3130 2502
rect 3086 2488 3090 2492
rect 3094 2488 3098 2492
rect 3110 2478 3114 2482
rect 3166 2478 3170 2482
rect 3078 2468 3082 2472
rect 3134 2468 3138 2472
rect 3158 2468 3162 2472
rect 3070 2448 3074 2452
rect 3142 2448 3146 2452
rect 3166 2448 3170 2452
rect 3118 2438 3122 2442
rect 3134 2438 3138 2442
rect 3094 2368 3098 2372
rect 3214 2658 3218 2662
rect 3198 2648 3202 2652
rect 3214 2648 3218 2652
rect 3182 2628 3186 2632
rect 3182 2618 3186 2622
rect 3230 2638 3234 2642
rect 3238 2638 3242 2642
rect 3550 2748 3554 2752
rect 3566 2738 3570 2742
rect 3582 2738 3586 2742
rect 3534 2718 3538 2722
rect 3526 2708 3530 2712
rect 3326 2658 3330 2662
rect 3414 2658 3418 2662
rect 3294 2648 3298 2652
rect 3262 2638 3266 2642
rect 3246 2628 3250 2632
rect 3246 2558 3250 2562
rect 3190 2538 3194 2542
rect 3238 2548 3242 2552
rect 3262 2548 3266 2552
rect 3206 2528 3210 2532
rect 3230 2538 3234 2542
rect 3310 2578 3314 2582
rect 3374 2628 3378 2632
rect 3342 2578 3346 2582
rect 3326 2568 3330 2572
rect 3326 2548 3330 2552
rect 3302 2538 3306 2542
rect 3342 2538 3346 2542
rect 3214 2518 3218 2522
rect 3214 2508 3218 2512
rect 3182 2488 3186 2492
rect 3198 2488 3202 2492
rect 3190 2478 3194 2482
rect 3254 2528 3258 2532
rect 3294 2528 3298 2532
rect 3334 2528 3338 2532
rect 3286 2518 3290 2522
rect 3318 2518 3322 2522
rect 3246 2498 3250 2502
rect 3278 2498 3282 2502
rect 3318 2498 3322 2502
rect 3222 2488 3226 2492
rect 3230 2488 3234 2492
rect 3318 2488 3322 2492
rect 3206 2468 3210 2472
rect 3254 2468 3258 2472
rect 3246 2458 3250 2462
rect 3270 2458 3274 2462
rect 3294 2468 3298 2472
rect 3318 2468 3322 2472
rect 3302 2458 3306 2462
rect 3358 2518 3362 2522
rect 3358 2488 3362 2492
rect 3542 2648 3546 2652
rect 3534 2638 3538 2642
rect 3518 2618 3522 2622
rect 3474 2603 3478 2607
rect 3481 2603 3485 2607
rect 3446 2598 3450 2602
rect 3462 2548 3466 2552
rect 3414 2498 3418 2502
rect 3486 2488 3490 2492
rect 3366 2468 3370 2472
rect 3382 2468 3386 2472
rect 3430 2468 3434 2472
rect 3446 2468 3450 2472
rect 3494 2478 3498 2482
rect 3494 2468 3498 2472
rect 3342 2458 3346 2462
rect 3358 2458 3362 2462
rect 3422 2458 3426 2462
rect 3278 2448 3282 2452
rect 3342 2448 3346 2452
rect 3174 2438 3178 2442
rect 3150 2428 3154 2432
rect 3166 2428 3170 2432
rect 3142 2418 3146 2422
rect 3166 2378 3170 2382
rect 3182 2378 3186 2382
rect 3262 2438 3266 2442
rect 3462 2448 3466 2452
rect 3398 2418 3402 2422
rect 3474 2403 3478 2407
rect 3481 2403 3485 2407
rect 3406 2388 3410 2392
rect 3238 2368 3242 2372
rect 3158 2358 3162 2362
rect 3190 2358 3194 2362
rect 3062 2348 3066 2352
rect 3174 2348 3178 2352
rect 3198 2348 3202 2352
rect 3222 2348 3226 2352
rect 3086 2338 3090 2342
rect 3134 2338 3138 2342
rect 3006 2328 3010 2332
rect 3070 2328 3074 2332
rect 3158 2328 3162 2332
rect 3078 2318 3082 2322
rect 3190 2308 3194 2312
rect 3134 2278 3138 2282
rect 3182 2278 3186 2282
rect 2998 2258 3002 2262
rect 3078 2258 3082 2262
rect 3030 2238 3034 2242
rect 3294 2358 3298 2362
rect 3326 2358 3330 2362
rect 3334 2358 3338 2362
rect 3470 2358 3474 2362
rect 3270 2348 3274 2352
rect 3302 2348 3306 2352
rect 3310 2348 3314 2352
rect 3254 2338 3258 2342
rect 3206 2328 3210 2332
rect 3214 2328 3218 2332
rect 3230 2328 3234 2332
rect 3206 2318 3210 2322
rect 3206 2298 3210 2302
rect 3198 2268 3202 2272
rect 3230 2318 3234 2322
rect 3278 2338 3282 2342
rect 3302 2338 3306 2342
rect 3358 2348 3362 2352
rect 3406 2348 3410 2352
rect 3342 2338 3346 2342
rect 3270 2328 3274 2332
rect 3278 2328 3282 2332
rect 3334 2328 3338 2332
rect 3262 2308 3266 2312
rect 3270 2308 3274 2312
rect 3302 2308 3306 2312
rect 3334 2318 3338 2322
rect 3358 2328 3362 2332
rect 3366 2318 3370 2322
rect 3342 2308 3346 2312
rect 3358 2298 3362 2302
rect 3398 2298 3402 2302
rect 3406 2298 3410 2302
rect 3326 2268 3330 2272
rect 3230 2258 3234 2262
rect 3118 2228 3122 2232
rect 2982 2198 2986 2202
rect 3078 2198 3082 2202
rect 2958 2188 2962 2192
rect 2910 2138 2914 2142
rect 2910 2128 2914 2132
rect 2806 2118 2810 2122
rect 2742 2108 2746 2112
rect 2750 2108 2754 2112
rect 2838 2108 2842 2112
rect 2894 2108 2898 2112
rect 2702 2088 2706 2092
rect 2734 2088 2738 2092
rect 2862 2098 2866 2102
rect 2774 2078 2778 2082
rect 2798 2078 2802 2082
rect 2830 2078 2834 2082
rect 2838 2078 2842 2082
rect 2718 2068 2722 2072
rect 2870 2088 2874 2092
rect 2902 2098 2906 2102
rect 2910 2088 2914 2092
rect 2990 2168 2994 2172
rect 2942 2138 2946 2142
rect 2954 2103 2958 2107
rect 2961 2103 2965 2107
rect 2926 2078 2930 2082
rect 2710 2058 2714 2062
rect 2846 2058 2850 2062
rect 2894 2058 2898 2062
rect 2918 2058 2922 2062
rect 2726 2048 2730 2052
rect 2758 2048 2762 2052
rect 2774 2048 2778 2052
rect 2750 2038 2754 2042
rect 2790 2038 2794 2042
rect 2806 2038 2810 2042
rect 2798 2028 2802 2032
rect 2742 2018 2746 2022
rect 2910 2038 2914 2042
rect 2822 2008 2826 2012
rect 2926 2008 2930 2012
rect 2846 1998 2850 2002
rect 2934 1998 2938 2002
rect 2950 1988 2954 1992
rect 2942 1968 2946 1972
rect 2766 1948 2770 1952
rect 2822 1948 2826 1952
rect 2886 1948 2890 1952
rect 2942 1948 2946 1952
rect 2974 1938 2978 1942
rect 2870 1928 2874 1932
rect 2750 1918 2754 1922
rect 2726 1908 2730 1912
rect 2718 1888 2722 1892
rect 2790 1898 2794 1902
rect 2694 1858 2698 1862
rect 2710 1858 2714 1862
rect 2734 1858 2738 1862
rect 2686 1848 2690 1852
rect 2718 1848 2722 1852
rect 2662 1818 2666 1822
rect 2606 1788 2610 1792
rect 2582 1758 2586 1762
rect 2654 1758 2658 1762
rect 2630 1748 2634 1752
rect 2558 1738 2562 1742
rect 2582 1738 2586 1742
rect 2606 1738 2610 1742
rect 2566 1718 2570 1722
rect 2574 1708 2578 1712
rect 2622 1718 2626 1722
rect 2590 1678 2594 1682
rect 2606 1658 2610 1662
rect 2630 1658 2634 1662
rect 2502 1648 2506 1652
rect 2606 1648 2610 1652
rect 2614 1648 2618 1652
rect 2638 1648 2642 1652
rect 2622 1628 2626 1632
rect 2442 1603 2446 1607
rect 2449 1603 2453 1607
rect 2534 1598 2538 1602
rect 2798 1858 2802 1862
rect 2806 1858 2810 1862
rect 2814 1858 2818 1862
rect 2878 1858 2882 1862
rect 2694 1838 2698 1842
rect 2742 1838 2746 1842
rect 2670 1728 2674 1732
rect 2686 1718 2690 1722
rect 2686 1688 2690 1692
rect 2654 1678 2658 1682
rect 2774 1838 2778 1842
rect 2750 1818 2754 1822
rect 2758 1818 2762 1822
rect 2710 1758 2714 1762
rect 2734 1758 2738 1762
rect 2798 1838 2802 1842
rect 2846 1818 2850 1822
rect 2878 1798 2882 1802
rect 2878 1778 2882 1782
rect 2814 1768 2818 1772
rect 2862 1768 2866 1772
rect 2758 1758 2762 1762
rect 2790 1758 2794 1762
rect 2822 1758 2826 1762
rect 2822 1748 2826 1752
rect 2766 1738 2770 1742
rect 2798 1738 2802 1742
rect 2710 1728 2714 1732
rect 2742 1728 2746 1732
rect 2774 1728 2778 1732
rect 2782 1728 2786 1732
rect 2702 1718 2706 1722
rect 2702 1698 2706 1702
rect 2758 1698 2762 1702
rect 2806 1698 2810 1702
rect 2750 1688 2754 1692
rect 2766 1688 2770 1692
rect 2782 1688 2786 1692
rect 2662 1638 2666 1642
rect 2646 1618 2650 1622
rect 2678 1618 2682 1622
rect 2678 1608 2682 1612
rect 2718 1658 2722 1662
rect 2710 1648 2714 1652
rect 2694 1598 2698 1602
rect 2718 1598 2722 1602
rect 2550 1558 2554 1562
rect 2606 1558 2610 1562
rect 2806 1678 2810 1682
rect 2758 1658 2762 1662
rect 2838 1728 2842 1732
rect 2870 1708 2874 1712
rect 2838 1698 2842 1702
rect 2862 1698 2866 1702
rect 2830 1688 2834 1692
rect 2918 1708 2922 1712
rect 2886 1688 2890 1692
rect 2846 1668 2850 1672
rect 2830 1638 2834 1642
rect 2846 1638 2850 1642
rect 2742 1628 2746 1632
rect 2734 1578 2738 1582
rect 2638 1558 2642 1562
rect 2686 1558 2690 1562
rect 2726 1558 2730 1562
rect 2734 1558 2738 1562
rect 2886 1558 2890 1562
rect 2438 1548 2442 1552
rect 2558 1548 2562 1552
rect 2574 1548 2578 1552
rect 2614 1548 2618 1552
rect 2654 1548 2658 1552
rect 2670 1548 2674 1552
rect 2422 1538 2426 1542
rect 2486 1528 2490 1532
rect 2526 1528 2530 1532
rect 2422 1518 2426 1522
rect 2510 1518 2514 1522
rect 2406 1488 2410 1492
rect 2510 1478 2514 1482
rect 2390 1468 2394 1472
rect 2454 1468 2458 1472
rect 2478 1468 2482 1472
rect 2590 1528 2594 1532
rect 2710 1548 2714 1552
rect 2638 1528 2642 1532
rect 2670 1528 2674 1532
rect 2598 1518 2602 1522
rect 2630 1518 2634 1522
rect 2558 1498 2562 1502
rect 2654 1498 2658 1502
rect 2686 1498 2690 1502
rect 2566 1488 2570 1492
rect 2782 1548 2786 1552
rect 2822 1548 2826 1552
rect 2886 1548 2890 1552
rect 2750 1538 2754 1542
rect 2782 1528 2786 1532
rect 2742 1518 2746 1522
rect 2718 1508 2722 1512
rect 2710 1488 2714 1492
rect 2694 1478 2698 1482
rect 2702 1478 2706 1482
rect 2734 1478 2738 1482
rect 2678 1468 2682 1472
rect 2422 1458 2426 1462
rect 2582 1458 2586 1462
rect 2638 1458 2642 1462
rect 2726 1468 2730 1472
rect 2398 1448 2402 1452
rect 2422 1448 2426 1452
rect 2478 1448 2482 1452
rect 2382 1418 2386 1422
rect 2438 1428 2442 1432
rect 2438 1418 2442 1422
rect 2510 1418 2514 1422
rect 2442 1403 2446 1407
rect 2449 1403 2453 1407
rect 2462 1398 2466 1402
rect 2438 1388 2442 1392
rect 2398 1358 2402 1362
rect 2390 1348 2394 1352
rect 2406 1348 2410 1352
rect 2102 1318 2106 1322
rect 2158 1318 2162 1322
rect 2198 1318 2202 1322
rect 2062 1288 2066 1292
rect 2206 1278 2210 1282
rect 2286 1278 2290 1282
rect 1990 1268 1994 1272
rect 2014 1268 2018 1272
rect 2030 1268 2034 1272
rect 2054 1268 2058 1272
rect 2070 1268 2074 1272
rect 2190 1268 2194 1272
rect 2006 1258 2010 1262
rect 1982 1248 1986 1252
rect 1966 1228 1970 1232
rect 1982 1158 1986 1162
rect 2062 1248 2066 1252
rect 2054 1218 2058 1222
rect 2102 1238 2106 1242
rect 2286 1258 2290 1262
rect 2278 1238 2282 1242
rect 2302 1238 2306 1242
rect 2318 1228 2322 1232
rect 2254 1218 2258 1222
rect 2150 1198 2154 1202
rect 2166 1198 2170 1202
rect 2174 1198 2178 1202
rect 2094 1188 2098 1192
rect 1982 1148 1986 1152
rect 2118 1148 2122 1152
rect 1950 1128 1954 1132
rect 1998 1128 2002 1132
rect 2014 1128 2018 1132
rect 1902 1118 1906 1122
rect 2014 1118 2018 1122
rect 2102 1118 2106 1122
rect 2150 1118 2154 1122
rect 1930 1103 1934 1107
rect 1937 1103 1941 1107
rect 2022 1108 2026 1112
rect 1950 1098 1954 1102
rect 2094 1098 2098 1102
rect 2118 1098 2122 1102
rect 1894 1088 1898 1092
rect 1918 1088 1922 1092
rect 1910 1078 1914 1082
rect 1966 1078 1970 1082
rect 1982 1078 1986 1082
rect 2022 1078 2026 1082
rect 2062 1078 2066 1082
rect 1926 1068 1930 1072
rect 2078 1068 2082 1072
rect 2102 1068 2106 1072
rect 1806 1038 1810 1042
rect 1782 1028 1786 1032
rect 1758 1018 1762 1022
rect 1822 1048 1826 1052
rect 1814 1008 1818 1012
rect 1774 978 1778 982
rect 1782 978 1786 982
rect 1758 958 1762 962
rect 1774 958 1778 962
rect 1758 938 1762 942
rect 1798 948 1802 952
rect 1854 1048 1858 1052
rect 1862 1008 1866 1012
rect 1846 958 1850 962
rect 1950 1058 1954 1062
rect 1910 1008 1914 1012
rect 1990 1038 1994 1042
rect 2030 1048 2034 1052
rect 1950 1018 1954 1022
rect 2006 1018 2010 1022
rect 2126 1078 2130 1082
rect 2094 1058 2098 1062
rect 2046 1008 2050 1012
rect 1998 978 2002 982
rect 2038 978 2042 982
rect 1878 958 1882 962
rect 1982 958 1986 962
rect 2054 958 2058 962
rect 1854 948 1858 952
rect 1878 948 1882 952
rect 1894 948 1898 952
rect 1926 948 1930 952
rect 1966 948 1970 952
rect 2038 948 2042 952
rect 2078 948 2082 952
rect 1790 938 1794 942
rect 1806 928 1810 932
rect 1758 878 1762 882
rect 1766 868 1770 872
rect 1782 878 1786 882
rect 1806 878 1810 882
rect 1830 938 1834 942
rect 1878 928 1882 932
rect 1830 878 1834 882
rect 1790 868 1794 872
rect 1814 868 1818 872
rect 1750 848 1754 852
rect 1798 838 1802 842
rect 1806 838 1810 842
rect 1806 828 1810 832
rect 1766 768 1770 772
rect 1782 758 1786 762
rect 1798 748 1802 752
rect 1846 868 1850 872
rect 1894 858 1898 862
rect 1870 848 1874 852
rect 1822 838 1826 842
rect 1926 928 1930 932
rect 2014 938 2018 942
rect 1958 918 1962 922
rect 1974 918 1978 922
rect 1930 903 1934 907
rect 1937 903 1941 907
rect 1982 888 1986 892
rect 1998 888 2002 892
rect 2126 1018 2130 1022
rect 2102 978 2106 982
rect 2198 1188 2202 1192
rect 2230 1158 2234 1162
rect 2374 1328 2378 1332
rect 2398 1328 2402 1332
rect 2430 1328 2434 1332
rect 2422 1278 2426 1282
rect 2406 1268 2410 1272
rect 2526 1398 2530 1402
rect 2566 1398 2570 1402
rect 2470 1388 2474 1392
rect 2510 1388 2514 1392
rect 2550 1388 2554 1392
rect 2478 1378 2482 1382
rect 2502 1378 2506 1382
rect 2486 1348 2490 1352
rect 2494 1348 2498 1352
rect 2526 1358 2530 1362
rect 2558 1378 2562 1382
rect 2614 1388 2618 1392
rect 2574 1358 2578 1362
rect 2582 1358 2586 1362
rect 2350 1208 2354 1212
rect 2442 1203 2446 1207
rect 2449 1203 2453 1207
rect 2302 1198 2306 1202
rect 2270 1168 2274 1172
rect 2430 1168 2434 1172
rect 2262 1158 2266 1162
rect 2318 1158 2322 1162
rect 2198 1148 2202 1152
rect 2214 1148 2218 1152
rect 2286 1148 2290 1152
rect 2302 1148 2306 1152
rect 2190 1118 2194 1122
rect 2206 1118 2210 1122
rect 2166 1078 2170 1082
rect 2142 1048 2146 1052
rect 2142 1008 2146 1012
rect 2134 968 2138 972
rect 2118 948 2122 952
rect 2286 1128 2290 1132
rect 2310 1128 2314 1132
rect 2342 1128 2346 1132
rect 2526 1328 2530 1332
rect 2518 1288 2522 1292
rect 2510 1258 2514 1262
rect 2486 1228 2490 1232
rect 2542 1258 2546 1262
rect 2598 1328 2602 1332
rect 2630 1378 2634 1382
rect 2622 1358 2626 1362
rect 2622 1318 2626 1322
rect 2654 1448 2658 1452
rect 2710 1418 2714 1422
rect 2954 1903 2958 1907
rect 2961 1903 2965 1907
rect 3254 2258 3258 2262
rect 3254 2248 3258 2252
rect 3246 2238 3250 2242
rect 3238 2228 3242 2232
rect 3230 2188 3234 2192
rect 3270 2188 3274 2192
rect 3262 2178 3266 2182
rect 3182 2168 3186 2172
rect 3238 2168 3242 2172
rect 3166 2148 3170 2152
rect 3094 2128 3098 2132
rect 3014 2078 3018 2082
rect 3102 2078 3106 2082
rect 2998 2058 3002 2062
rect 3006 1978 3010 1982
rect 3198 2148 3202 2152
rect 3246 2148 3250 2152
rect 3278 2178 3282 2182
rect 3294 2248 3298 2252
rect 3302 2218 3306 2222
rect 3318 2238 3322 2242
rect 3326 2238 3330 2242
rect 3526 2478 3530 2482
rect 3590 2718 3594 2722
rect 3614 2848 3618 2852
rect 3654 2858 3658 2862
rect 3678 2848 3682 2852
rect 3630 2828 3634 2832
rect 3646 2808 3650 2812
rect 3670 2838 3674 2842
rect 3654 2768 3658 2772
rect 3710 2908 3714 2912
rect 3718 2898 3722 2902
rect 3710 2888 3714 2892
rect 3758 2928 3762 2932
rect 3926 3068 3930 3072
rect 3974 3068 3978 3072
rect 4038 3068 4042 3072
rect 4086 3068 4090 3072
rect 4142 3068 4146 3072
rect 3878 3058 3882 3062
rect 3902 3058 3906 3062
rect 3862 3038 3866 3042
rect 3894 3038 3898 3042
rect 3886 3018 3890 3022
rect 3878 2998 3882 3002
rect 3854 2978 3858 2982
rect 3934 3048 3938 3052
rect 3950 3048 3954 3052
rect 3910 3018 3914 3022
rect 3958 3018 3962 3022
rect 3902 2998 3906 3002
rect 3958 2998 3962 3002
rect 3894 2958 3898 2962
rect 3950 2958 3954 2962
rect 3958 2958 3962 2962
rect 3838 2928 3842 2932
rect 3926 2928 3930 2932
rect 3766 2888 3770 2892
rect 3790 2888 3794 2892
rect 3702 2868 3706 2872
rect 3782 2868 3786 2872
rect 3774 2858 3778 2862
rect 3806 2858 3810 2862
rect 3926 2918 3930 2922
rect 3886 2888 3890 2892
rect 3862 2868 3866 2872
rect 3886 2868 3890 2872
rect 3910 2868 3914 2872
rect 3838 2858 3842 2862
rect 3894 2858 3898 2862
rect 3798 2848 3802 2852
rect 3814 2848 3818 2852
rect 3854 2848 3858 2852
rect 3838 2838 3842 2842
rect 3886 2838 3890 2842
rect 3910 2838 3914 2842
rect 3838 2828 3842 2832
rect 3854 2828 3858 2832
rect 3878 2828 3882 2832
rect 3702 2818 3706 2822
rect 3742 2808 3746 2812
rect 3774 2808 3778 2812
rect 3814 2808 3818 2812
rect 3662 2758 3666 2762
rect 3646 2748 3650 2752
rect 3750 2748 3754 2752
rect 3646 2728 3650 2732
rect 3598 2708 3602 2712
rect 3606 2708 3610 2712
rect 3582 2698 3586 2702
rect 3582 2688 3586 2692
rect 3566 2678 3570 2682
rect 3582 2668 3586 2672
rect 3614 2688 3618 2692
rect 3614 2668 3618 2672
rect 3558 2658 3562 2662
rect 3574 2648 3578 2652
rect 3550 2628 3554 2632
rect 3790 2768 3794 2772
rect 3782 2748 3786 2752
rect 3798 2748 3802 2752
rect 3806 2748 3810 2752
rect 3718 2728 3722 2732
rect 3734 2728 3738 2732
rect 3758 2728 3762 2732
rect 3654 2718 3658 2722
rect 3694 2718 3698 2722
rect 3678 2698 3682 2702
rect 3710 2698 3714 2702
rect 3702 2688 3706 2692
rect 3806 2688 3810 2692
rect 3774 2678 3778 2682
rect 3790 2678 3794 2682
rect 3998 3058 4002 3062
rect 4006 3058 4010 3062
rect 4022 3058 4026 3062
rect 4062 3058 4066 3062
rect 4102 3058 4106 3062
rect 4110 3058 4114 3062
rect 3998 3048 4002 3052
rect 3982 2948 3986 2952
rect 4038 3048 4042 3052
rect 4030 3038 4034 3042
rect 4110 3038 4114 3042
rect 4102 3028 4106 3032
rect 4126 3028 4130 3032
rect 4054 3008 4058 3012
rect 4046 2998 4050 3002
rect 4102 2988 4106 2992
rect 3998 2978 4002 2982
rect 4054 2978 4058 2982
rect 4110 2978 4114 2982
rect 4038 2968 4042 2972
rect 4022 2948 4026 2952
rect 3990 2918 3994 2922
rect 3978 2903 3982 2907
rect 3985 2903 3989 2907
rect 3998 2898 4002 2902
rect 3934 2888 3938 2892
rect 3966 2888 3970 2892
rect 4198 3068 4202 3072
rect 4238 3068 4242 3072
rect 4254 3068 4258 3072
rect 4286 3068 4290 3072
rect 4302 3058 4306 3062
rect 4158 3048 4162 3052
rect 4174 3038 4178 3042
rect 4166 3018 4170 3022
rect 4142 3008 4146 3012
rect 4190 3028 4194 3032
rect 4198 2978 4202 2982
rect 4086 2968 4090 2972
rect 4118 2968 4122 2972
rect 4134 2968 4138 2972
rect 4150 2968 4154 2972
rect 4166 2968 4170 2972
rect 4182 2968 4186 2972
rect 4014 2928 4018 2932
rect 4046 2928 4050 2932
rect 4094 2958 4098 2962
rect 4150 2958 4154 2962
rect 4174 2958 4178 2962
rect 4118 2948 4122 2952
rect 4158 2948 4162 2952
rect 4070 2938 4074 2942
rect 4102 2938 4106 2942
rect 4086 2928 4090 2932
rect 4150 2928 4154 2932
rect 4030 2908 4034 2912
rect 4062 2908 4066 2912
rect 4134 2908 4138 2912
rect 4190 2948 4194 2952
rect 4214 2988 4218 2992
rect 4198 2928 4202 2932
rect 4206 2928 4210 2932
rect 4270 3048 4274 3052
rect 4294 3048 4298 3052
rect 4310 3038 4314 3042
rect 4246 3028 4250 3032
rect 4294 3028 4298 3032
rect 4238 3018 4242 3022
rect 4238 2998 4242 3002
rect 4294 3008 4298 3012
rect 4262 2998 4266 3002
rect 4342 2998 4346 3002
rect 4374 2988 4378 2992
rect 4374 2978 4378 2982
rect 4262 2968 4266 2972
rect 4326 2968 4330 2972
rect 4254 2948 4258 2952
rect 4230 2928 4234 2932
rect 4222 2918 4226 2922
rect 4238 2918 4242 2922
rect 4254 2918 4258 2922
rect 4182 2908 4186 2912
rect 4166 2898 4170 2902
rect 4174 2898 4178 2902
rect 4230 2908 4234 2912
rect 4030 2888 4034 2892
rect 4038 2888 4042 2892
rect 4206 2888 4210 2892
rect 3982 2878 3986 2882
rect 3942 2868 3946 2872
rect 3958 2868 3962 2872
rect 3926 2858 3930 2862
rect 3966 2858 3970 2862
rect 3950 2848 3954 2852
rect 3974 2848 3978 2852
rect 3934 2828 3938 2832
rect 3918 2808 3922 2812
rect 3886 2778 3890 2782
rect 3878 2768 3882 2772
rect 3846 2748 3850 2752
rect 3870 2748 3874 2752
rect 3838 2738 3842 2742
rect 3838 2728 3842 2732
rect 3942 2758 3946 2762
rect 3894 2748 3898 2752
rect 3982 2748 3986 2752
rect 3870 2728 3874 2732
rect 3854 2718 3858 2722
rect 3822 2678 3826 2682
rect 3934 2728 3938 2732
rect 3902 2708 3906 2712
rect 3766 2668 3770 2672
rect 3734 2658 3738 2662
rect 3774 2658 3778 2662
rect 3606 2618 3610 2622
rect 3630 2618 3634 2622
rect 3638 2608 3642 2612
rect 3670 2648 3674 2652
rect 3734 2648 3738 2652
rect 3766 2618 3770 2622
rect 3694 2598 3698 2602
rect 3558 2578 3562 2582
rect 3662 2578 3666 2582
rect 3550 2528 3554 2532
rect 3534 2468 3538 2472
rect 3542 2468 3546 2472
rect 3630 2558 3634 2562
rect 3646 2558 3650 2562
rect 3694 2558 3698 2562
rect 3590 2548 3594 2552
rect 3614 2538 3618 2542
rect 3606 2528 3610 2532
rect 3566 2518 3570 2522
rect 3614 2518 3618 2522
rect 3566 2508 3570 2512
rect 3590 2488 3594 2492
rect 3614 2478 3618 2482
rect 3622 2468 3626 2472
rect 3838 2668 3842 2672
rect 3886 2678 3890 2682
rect 3894 2668 3898 2672
rect 3870 2658 3874 2662
rect 3854 2638 3858 2642
rect 3838 2628 3842 2632
rect 3790 2618 3794 2622
rect 3846 2608 3850 2612
rect 3918 2678 3922 2682
rect 3910 2648 3914 2652
rect 3902 2628 3906 2632
rect 3854 2598 3858 2602
rect 3814 2558 3818 2562
rect 3774 2548 3778 2552
rect 3782 2548 3786 2552
rect 3806 2548 3810 2552
rect 3654 2528 3658 2532
rect 3686 2538 3690 2542
rect 3710 2538 3714 2542
rect 3766 2538 3770 2542
rect 3670 2528 3674 2532
rect 3662 2498 3666 2502
rect 3726 2508 3730 2512
rect 3662 2488 3666 2492
rect 3694 2488 3698 2492
rect 3654 2478 3658 2482
rect 3710 2478 3714 2482
rect 3686 2468 3690 2472
rect 3718 2468 3722 2472
rect 3758 2528 3762 2532
rect 3774 2528 3778 2532
rect 3774 2508 3778 2512
rect 3742 2498 3746 2502
rect 3782 2488 3786 2492
rect 3830 2538 3834 2542
rect 3846 2538 3850 2542
rect 3526 2458 3530 2462
rect 3630 2458 3634 2462
rect 3662 2458 3666 2462
rect 3774 2458 3778 2462
rect 3814 2458 3818 2462
rect 3542 2448 3546 2452
rect 3550 2368 3554 2372
rect 3518 2348 3522 2352
rect 3502 2318 3506 2322
rect 3454 2288 3458 2292
rect 3414 2278 3418 2282
rect 3430 2278 3434 2282
rect 3502 2278 3506 2282
rect 3422 2268 3426 2272
rect 3462 2268 3466 2272
rect 3374 2258 3378 2262
rect 3390 2258 3394 2262
rect 3406 2258 3410 2262
rect 3454 2258 3458 2262
rect 3350 2248 3354 2252
rect 3382 2248 3386 2252
rect 3478 2248 3482 2252
rect 3486 2248 3490 2252
rect 3454 2228 3458 2232
rect 3334 2208 3338 2212
rect 3494 2208 3498 2212
rect 3474 2203 3478 2207
rect 3481 2203 3485 2207
rect 3374 2178 3378 2182
rect 3414 2178 3418 2182
rect 3422 2178 3426 2182
rect 3470 2168 3474 2172
rect 3286 2158 3290 2162
rect 3566 2448 3570 2452
rect 3558 2338 3562 2342
rect 3606 2428 3610 2432
rect 3654 2428 3658 2432
rect 3798 2428 3802 2432
rect 3630 2378 3634 2382
rect 3582 2368 3586 2372
rect 3838 2518 3842 2522
rect 3886 2588 3890 2592
rect 3934 2658 3938 2662
rect 3926 2648 3930 2652
rect 3966 2728 3970 2732
rect 3974 2728 3978 2732
rect 3950 2658 3954 2662
rect 3982 2718 3986 2722
rect 3978 2703 3982 2707
rect 3985 2703 3989 2707
rect 4006 2878 4010 2882
rect 4006 2868 4010 2872
rect 4030 2868 4034 2872
rect 4014 2858 4018 2862
rect 4006 2778 4010 2782
rect 3998 2688 4002 2692
rect 3982 2678 3986 2682
rect 3958 2648 3962 2652
rect 4006 2648 4010 2652
rect 3934 2628 3938 2632
rect 3950 2628 3954 2632
rect 3918 2548 3922 2552
rect 3966 2598 3970 2602
rect 4006 2588 4010 2592
rect 3974 2558 3978 2562
rect 3950 2538 3954 2542
rect 4246 2878 4250 2882
rect 4062 2868 4066 2872
rect 4094 2868 4098 2872
rect 4126 2868 4130 2872
rect 4134 2868 4138 2872
rect 4214 2868 4218 2872
rect 4246 2868 4250 2872
rect 4054 2858 4058 2862
rect 4086 2858 4090 2862
rect 4118 2858 4122 2862
rect 4046 2838 4050 2842
rect 4078 2818 4082 2822
rect 4038 2798 4042 2802
rect 4030 2788 4034 2792
rect 4062 2748 4066 2752
rect 4070 2738 4074 2742
rect 4038 2728 4042 2732
rect 4078 2718 4082 2722
rect 4054 2708 4058 2712
rect 4030 2688 4034 2692
rect 4046 2678 4050 2682
rect 4142 2858 4146 2862
rect 4198 2858 4202 2862
rect 4214 2858 4218 2862
rect 4334 2958 4338 2962
rect 4342 2958 4346 2962
rect 4366 2958 4370 2962
rect 4310 2948 4314 2952
rect 4318 2948 4322 2952
rect 4286 2918 4290 2922
rect 4294 2898 4298 2902
rect 4278 2878 4282 2882
rect 4286 2878 4290 2882
rect 4270 2868 4274 2872
rect 4126 2788 4130 2792
rect 4110 2768 4114 2772
rect 4118 2728 4122 2732
rect 4134 2728 4138 2732
rect 4030 2668 4034 2672
rect 4102 2668 4106 2672
rect 4126 2718 4130 2722
rect 4182 2818 4186 2822
rect 4150 2788 4154 2792
rect 4278 2848 4282 2852
rect 4206 2808 4210 2812
rect 4246 2808 4250 2812
rect 4222 2798 4226 2802
rect 4190 2778 4194 2782
rect 4214 2778 4218 2782
rect 4182 2748 4186 2752
rect 4166 2738 4170 2742
rect 4182 2698 4186 2702
rect 4198 2758 4202 2762
rect 4198 2748 4202 2752
rect 4246 2748 4250 2752
rect 4270 2748 4274 2752
rect 4142 2678 4146 2682
rect 4174 2678 4178 2682
rect 4046 2648 4050 2652
rect 4110 2648 4114 2652
rect 4022 2628 4026 2632
rect 4038 2588 4042 2592
rect 4014 2578 4018 2582
rect 4014 2538 4018 2542
rect 3870 2528 3874 2532
rect 3942 2528 3946 2532
rect 3966 2528 3970 2532
rect 3998 2528 4002 2532
rect 3894 2508 3898 2512
rect 3862 2488 3866 2492
rect 3894 2488 3898 2492
rect 3918 2478 3922 2482
rect 3862 2468 3866 2472
rect 3950 2518 3954 2522
rect 3978 2503 3982 2507
rect 3985 2503 3989 2507
rect 3966 2488 3970 2492
rect 3982 2488 3986 2492
rect 3934 2458 3938 2462
rect 3982 2458 3986 2462
rect 4030 2538 4034 2542
rect 4134 2658 4138 2662
rect 4142 2648 4146 2652
rect 4166 2648 4170 2652
rect 4126 2638 4130 2642
rect 4158 2638 4162 2642
rect 4118 2628 4122 2632
rect 4158 2628 4162 2632
rect 4078 2608 4082 2612
rect 4150 2598 4154 2602
rect 4142 2588 4146 2592
rect 4078 2568 4082 2572
rect 4054 2558 4058 2562
rect 4062 2558 4066 2562
rect 4070 2548 4074 2552
rect 4022 2528 4026 2532
rect 4062 2528 4066 2532
rect 4022 2478 4026 2482
rect 4134 2548 4138 2552
rect 4142 2538 4146 2542
rect 4126 2528 4130 2532
rect 4086 2518 4090 2522
rect 4078 2478 4082 2482
rect 4078 2468 4082 2472
rect 4070 2458 4074 2462
rect 4086 2458 4090 2462
rect 4022 2448 4026 2452
rect 3846 2438 3850 2442
rect 3926 2438 3930 2442
rect 3998 2438 4002 2442
rect 4094 2438 4098 2442
rect 3998 2428 4002 2432
rect 3822 2378 3826 2382
rect 3798 2368 3802 2372
rect 3582 2358 3586 2362
rect 3598 2358 3602 2362
rect 3574 2338 3578 2342
rect 3630 2348 3634 2352
rect 3822 2358 3826 2362
rect 3902 2368 3906 2372
rect 3926 2368 3930 2372
rect 3846 2358 3850 2362
rect 3894 2358 3898 2362
rect 3902 2358 3906 2362
rect 4054 2368 4058 2372
rect 4006 2348 4010 2352
rect 4014 2348 4018 2352
rect 3814 2338 3818 2342
rect 3862 2338 3866 2342
rect 3622 2328 3626 2332
rect 3590 2318 3594 2322
rect 3614 2318 3618 2322
rect 3590 2298 3594 2302
rect 3606 2288 3610 2292
rect 3854 2328 3858 2332
rect 3678 2288 3682 2292
rect 3542 2268 3546 2272
rect 3550 2258 3554 2262
rect 3566 2258 3570 2262
rect 3582 2258 3586 2262
rect 3590 2258 3594 2262
rect 3526 2248 3530 2252
rect 3558 2248 3562 2252
rect 3526 2228 3530 2232
rect 3518 2188 3522 2192
rect 3526 2168 3530 2172
rect 3542 2168 3546 2172
rect 3510 2158 3514 2162
rect 3286 2148 3290 2152
rect 3350 2148 3354 2152
rect 3414 2148 3418 2152
rect 3238 2138 3242 2142
rect 3254 2138 3258 2142
rect 3206 2128 3210 2132
rect 3278 2128 3282 2132
rect 3214 2108 3218 2112
rect 3206 2098 3210 2102
rect 3166 2088 3170 2092
rect 3198 2088 3202 2092
rect 3182 2078 3186 2082
rect 3230 2088 3234 2092
rect 3254 2088 3258 2092
rect 3270 2088 3274 2092
rect 3214 2078 3218 2082
rect 3246 2078 3250 2082
rect 3254 2078 3258 2082
rect 3190 2068 3194 2072
rect 3198 2068 3202 2072
rect 3230 2068 3234 2072
rect 3198 2058 3202 2062
rect 3206 2058 3210 2062
rect 3086 2048 3090 2052
rect 3166 2048 3170 2052
rect 3134 2038 3138 2042
rect 3086 2018 3090 2022
rect 3054 2008 3058 2012
rect 3062 1968 3066 1972
rect 2998 1948 3002 1952
rect 3046 1948 3050 1952
rect 3094 1978 3098 1982
rect 3070 1958 3074 1962
rect 3182 1998 3186 2002
rect 3110 1958 3114 1962
rect 3166 1958 3170 1962
rect 3126 1948 3130 1952
rect 3142 1948 3146 1952
rect 3022 1938 3026 1942
rect 3086 1938 3090 1942
rect 3062 1928 3066 1932
rect 3094 1928 3098 1932
rect 3118 1938 3122 1942
rect 3062 1918 3066 1922
rect 3102 1918 3106 1922
rect 2982 1898 2986 1902
rect 3246 2038 3250 2042
rect 3230 2028 3234 2032
rect 3214 1978 3218 1982
rect 3206 1958 3210 1962
rect 3318 2138 3322 2142
rect 3342 2138 3346 2142
rect 3310 2098 3314 2102
rect 3302 2088 3306 2092
rect 3278 2078 3282 2082
rect 3262 2048 3266 2052
rect 3278 2048 3282 2052
rect 3310 2058 3314 2062
rect 3286 1998 3290 2002
rect 3294 1998 3298 2002
rect 3310 1998 3314 2002
rect 3286 1978 3290 1982
rect 3198 1948 3202 1952
rect 3222 1948 3226 1952
rect 3174 1938 3178 1942
rect 3254 1938 3258 1942
rect 3270 1938 3274 1942
rect 3310 1938 3314 1942
rect 3158 1928 3162 1932
rect 3206 1928 3210 1932
rect 3254 1928 3258 1932
rect 3126 1918 3130 1922
rect 3182 1918 3186 1922
rect 3118 1898 3122 1902
rect 3142 1898 3146 1902
rect 3174 1898 3178 1902
rect 3110 1888 3114 1892
rect 2950 1878 2954 1882
rect 2998 1878 3002 1882
rect 2942 1858 2946 1862
rect 2974 1858 2978 1862
rect 3126 1888 3130 1892
rect 3158 1888 3162 1892
rect 3086 1868 3090 1872
rect 3102 1868 3106 1872
rect 3078 1858 3082 1862
rect 3038 1818 3042 1822
rect 3078 1848 3082 1852
rect 3086 1848 3090 1852
rect 3214 1888 3218 1892
rect 3182 1868 3186 1872
rect 3198 1868 3202 1872
rect 3238 1868 3242 1872
rect 3326 2128 3330 2132
rect 3374 2138 3378 2142
rect 3358 2118 3362 2122
rect 3422 2138 3426 2142
rect 3462 2138 3466 2142
rect 3414 2128 3418 2132
rect 3446 2128 3450 2132
rect 3462 2128 3466 2132
rect 3390 2118 3394 2122
rect 3358 2108 3362 2112
rect 3382 2108 3386 2112
rect 3334 2098 3338 2102
rect 3382 2088 3386 2092
rect 3438 2108 3442 2112
rect 3406 2078 3410 2082
rect 3422 2078 3426 2082
rect 3326 2068 3330 2072
rect 3342 2068 3346 2072
rect 3326 2058 3330 2062
rect 3326 2048 3330 2052
rect 3342 2038 3346 2042
rect 3374 2068 3378 2072
rect 3406 2068 3410 2072
rect 3502 2108 3506 2112
rect 3462 2098 3466 2102
rect 3494 2088 3498 2092
rect 3454 2078 3458 2082
rect 3470 2078 3474 2082
rect 3454 2058 3458 2062
rect 3366 2048 3370 2052
rect 3390 2018 3394 2022
rect 3358 1998 3362 2002
rect 3406 2048 3410 2052
rect 3398 1988 3402 1992
rect 3414 1978 3418 1982
rect 3406 1958 3410 1962
rect 3350 1948 3354 1952
rect 3430 1968 3434 1972
rect 3422 1958 3426 1962
rect 3438 1948 3442 1952
rect 3446 1948 3450 1952
rect 3542 2138 3546 2142
rect 3542 2088 3546 2092
rect 3518 2078 3522 2082
rect 3526 2068 3530 2072
rect 3550 2058 3554 2062
rect 3574 2248 3578 2252
rect 3606 2238 3610 2242
rect 3566 2228 3570 2232
rect 3606 2198 3610 2202
rect 3590 2178 3594 2182
rect 3590 2168 3594 2172
rect 3566 2158 3570 2162
rect 3566 2118 3570 2122
rect 3582 2128 3586 2132
rect 3574 2088 3578 2092
rect 3486 2048 3490 2052
rect 3518 2038 3522 2042
rect 3526 2038 3530 2042
rect 3474 2003 3478 2007
rect 3481 2003 3485 2007
rect 3510 1968 3514 1972
rect 3526 1988 3530 1992
rect 3694 2278 3698 2282
rect 4006 2328 4010 2332
rect 3894 2318 3898 2322
rect 3934 2318 3938 2322
rect 3950 2318 3954 2322
rect 3766 2308 3770 2312
rect 3662 2268 3666 2272
rect 3646 2258 3650 2262
rect 3630 2248 3634 2252
rect 3654 2248 3658 2252
rect 3662 2228 3666 2232
rect 3638 2148 3642 2152
rect 3614 2128 3618 2132
rect 3638 2108 3642 2112
rect 3622 2068 3626 2072
rect 3638 2068 3642 2072
rect 3590 2048 3594 2052
rect 3638 2058 3642 2062
rect 3574 2038 3578 2042
rect 3606 2038 3610 2042
rect 3598 2018 3602 2022
rect 3582 2008 3586 2012
rect 3542 1958 3546 1962
rect 3558 1958 3562 1962
rect 3534 1948 3538 1952
rect 3558 1948 3562 1952
rect 3358 1938 3362 1942
rect 3406 1938 3410 1942
rect 3462 1938 3466 1942
rect 3286 1928 3290 1932
rect 3318 1928 3322 1932
rect 3278 1918 3282 1922
rect 3398 1928 3402 1932
rect 3438 1918 3442 1922
rect 3350 1908 3354 1912
rect 3294 1898 3298 1902
rect 3150 1858 3154 1862
rect 3174 1858 3178 1862
rect 3206 1858 3210 1862
rect 3246 1858 3250 1862
rect 3190 1848 3194 1852
rect 3118 1818 3122 1822
rect 3142 1818 3146 1822
rect 3046 1798 3050 1802
rect 3014 1758 3018 1762
rect 3214 1778 3218 1782
rect 3102 1758 3106 1762
rect 3142 1758 3146 1762
rect 3174 1758 3178 1762
rect 3182 1758 3186 1762
rect 3086 1748 3090 1752
rect 3126 1748 3130 1752
rect 3166 1748 3170 1752
rect 3190 1748 3194 1752
rect 3118 1738 3122 1742
rect 3150 1738 3154 1742
rect 2998 1708 3002 1712
rect 3030 1708 3034 1712
rect 3054 1708 3058 1712
rect 2954 1703 2958 1707
rect 2961 1703 2965 1707
rect 2974 1698 2978 1702
rect 3142 1728 3146 1732
rect 3166 1718 3170 1722
rect 3086 1708 3090 1712
rect 3078 1698 3082 1702
rect 3190 1708 3194 1712
rect 3198 1708 3202 1712
rect 3174 1698 3178 1702
rect 3070 1668 3074 1672
rect 3158 1658 3162 1662
rect 3206 1658 3210 1662
rect 3134 1648 3138 1652
rect 3126 1628 3130 1632
rect 2966 1618 2970 1622
rect 2982 1618 2986 1622
rect 2942 1548 2946 1552
rect 2982 1548 2986 1552
rect 2982 1518 2986 1522
rect 2870 1508 2874 1512
rect 2910 1508 2914 1512
rect 2926 1508 2930 1512
rect 2774 1488 2778 1492
rect 2798 1488 2802 1492
rect 2750 1468 2754 1472
rect 2782 1468 2786 1472
rect 2838 1478 2842 1482
rect 2806 1468 2810 1472
rect 2846 1468 2850 1472
rect 2734 1448 2738 1452
rect 2750 1448 2754 1452
rect 2766 1448 2770 1452
rect 2734 1418 2738 1422
rect 2670 1408 2674 1412
rect 2718 1408 2722 1412
rect 2662 1358 2666 1362
rect 2654 1348 2658 1352
rect 2726 1378 2730 1382
rect 2686 1358 2690 1362
rect 2830 1458 2834 1462
rect 2790 1448 2794 1452
rect 2814 1428 2818 1432
rect 2838 1428 2842 1432
rect 2878 1458 2882 1462
rect 2894 1458 2898 1462
rect 2854 1418 2858 1422
rect 2846 1398 2850 1402
rect 2790 1368 2794 1372
rect 2814 1368 2818 1372
rect 2830 1368 2834 1372
rect 2806 1358 2810 1362
rect 2886 1408 2890 1412
rect 2686 1348 2690 1352
rect 2718 1348 2722 1352
rect 2774 1348 2778 1352
rect 2806 1348 2810 1352
rect 2742 1338 2746 1342
rect 2654 1328 2658 1332
rect 2710 1328 2714 1332
rect 2750 1328 2754 1332
rect 2798 1338 2802 1342
rect 2814 1338 2818 1342
rect 2862 1338 2866 1342
rect 2638 1308 2642 1312
rect 2670 1308 2674 1312
rect 2630 1288 2634 1292
rect 2694 1278 2698 1282
rect 2726 1288 2730 1292
rect 2742 1278 2746 1282
rect 2702 1268 2706 1272
rect 2734 1268 2738 1272
rect 2766 1268 2770 1272
rect 2574 1228 2578 1232
rect 2558 1218 2562 1222
rect 2606 1218 2610 1222
rect 2566 1158 2570 1162
rect 2582 1158 2586 1162
rect 2526 1148 2530 1152
rect 2550 1148 2554 1152
rect 2526 1128 2530 1132
rect 2238 1118 2242 1122
rect 2246 1118 2250 1122
rect 2318 1118 2322 1122
rect 2390 1118 2394 1122
rect 2446 1118 2450 1122
rect 2294 1098 2298 1102
rect 2222 1078 2226 1082
rect 2262 1068 2266 1072
rect 2350 1108 2354 1112
rect 2398 1108 2402 1112
rect 2438 1108 2442 1112
rect 2342 1098 2346 1102
rect 2326 1078 2330 1082
rect 2278 1048 2282 1052
rect 2382 1088 2386 1092
rect 2390 1058 2394 1062
rect 2350 1048 2354 1052
rect 2214 1008 2218 1012
rect 2326 1008 2330 1012
rect 2342 1008 2346 1012
rect 2238 978 2242 982
rect 2182 968 2186 972
rect 2094 918 2098 922
rect 2150 938 2154 942
rect 2166 938 2170 942
rect 2198 938 2202 942
rect 2118 928 2122 932
rect 2134 928 2138 932
rect 2150 928 2154 932
rect 2094 878 2098 882
rect 1982 868 1986 872
rect 2054 868 2058 872
rect 1942 848 1946 852
rect 1934 838 1938 842
rect 1910 828 1914 832
rect 1862 778 1866 782
rect 1854 748 1858 752
rect 1766 738 1770 742
rect 1774 688 1778 692
rect 1806 738 1810 742
rect 1814 708 1818 712
rect 1790 688 1794 692
rect 1750 678 1754 682
rect 1782 678 1786 682
rect 1734 658 1738 662
rect 1742 658 1746 662
rect 1758 658 1762 662
rect 1790 658 1794 662
rect 1718 648 1722 652
rect 1726 648 1730 652
rect 1686 638 1690 642
rect 1694 638 1698 642
rect 1678 578 1682 582
rect 1742 638 1746 642
rect 1694 568 1698 572
rect 1710 568 1714 572
rect 1742 558 1746 562
rect 1686 548 1690 552
rect 1766 638 1770 642
rect 1782 568 1786 572
rect 1798 568 1802 572
rect 1838 718 1842 722
rect 1846 698 1850 702
rect 1822 688 1826 692
rect 1822 678 1826 682
rect 1790 558 1794 562
rect 1806 558 1810 562
rect 1774 548 1778 552
rect 1670 538 1674 542
rect 1638 488 1642 492
rect 1614 458 1618 462
rect 1566 448 1570 452
rect 1582 428 1586 432
rect 1574 378 1578 382
rect 1566 368 1570 372
rect 1558 348 1562 352
rect 1566 348 1570 352
rect 1606 408 1610 412
rect 1590 358 1594 362
rect 1590 338 1594 342
rect 1566 318 1570 322
rect 1558 288 1562 292
rect 1598 308 1602 312
rect 1574 268 1578 272
rect 1462 258 1466 262
rect 1470 258 1474 262
rect 1502 258 1506 262
rect 1550 258 1554 262
rect 1478 248 1482 252
rect 1526 248 1530 252
rect 1454 228 1458 232
rect 1446 198 1450 202
rect 1470 228 1474 232
rect 1462 188 1466 192
rect 1454 158 1458 162
rect 1486 218 1490 222
rect 1494 178 1498 182
rect 1550 228 1554 232
rect 1494 158 1498 162
rect 1518 158 1522 162
rect 1534 158 1538 162
rect 1398 148 1402 152
rect 1414 148 1418 152
rect 1526 148 1530 152
rect 1566 218 1570 222
rect 1558 148 1562 152
rect 1454 138 1458 142
rect 1534 138 1538 142
rect 1614 278 1618 282
rect 1622 278 1626 282
rect 1590 248 1594 252
rect 1582 198 1586 202
rect 1590 178 1594 182
rect 1590 158 1594 162
rect 1598 158 1602 162
rect 1614 238 1618 242
rect 1654 478 1658 482
rect 1710 538 1714 542
rect 1726 538 1730 542
rect 1814 548 1818 552
rect 1814 538 1818 542
rect 1750 528 1754 532
rect 1774 528 1778 532
rect 1806 528 1810 532
rect 1750 488 1754 492
rect 1766 488 1770 492
rect 1710 478 1714 482
rect 1790 478 1794 482
rect 1654 448 1658 452
rect 1646 438 1650 442
rect 1646 418 1650 422
rect 1638 278 1642 282
rect 1670 398 1674 402
rect 1742 458 1746 462
rect 1766 458 1770 462
rect 1782 458 1786 462
rect 1774 448 1778 452
rect 1798 448 1802 452
rect 1734 438 1738 442
rect 1710 378 1714 382
rect 1694 368 1698 372
rect 1750 338 1754 342
rect 1694 328 1698 332
rect 1710 328 1714 332
rect 1670 288 1674 292
rect 1726 288 1730 292
rect 1822 518 1826 522
rect 1830 488 1834 492
rect 1822 478 1826 482
rect 1846 568 1850 572
rect 1886 758 1890 762
rect 1950 808 1954 812
rect 2046 838 2050 842
rect 2070 838 2074 842
rect 2078 798 2082 802
rect 2014 768 2018 772
rect 2038 758 2042 762
rect 2070 758 2074 762
rect 1926 748 1930 752
rect 1974 748 1978 752
rect 2022 748 2026 752
rect 2038 748 2042 752
rect 1894 728 1898 732
rect 1918 728 1922 732
rect 1870 708 1874 712
rect 1910 708 1914 712
rect 1902 688 1906 692
rect 1886 678 1890 682
rect 1894 658 1898 662
rect 1870 548 1874 552
rect 1974 708 1978 712
rect 1930 703 1934 707
rect 1937 703 1941 707
rect 1942 668 1946 672
rect 1910 588 1914 592
rect 1918 588 1922 592
rect 1910 578 1914 582
rect 1894 548 1898 552
rect 1854 538 1858 542
rect 1878 538 1882 542
rect 1854 528 1858 532
rect 1814 470 1818 472
rect 1814 468 1818 470
rect 1838 468 1842 472
rect 1862 458 1866 462
rect 1830 448 1834 452
rect 1806 318 1810 322
rect 1782 278 1786 282
rect 1798 278 1802 282
rect 1822 308 1826 312
rect 1814 298 1818 302
rect 1862 448 1866 452
rect 1854 408 1858 412
rect 1838 398 1842 402
rect 1838 378 1842 382
rect 1854 358 1858 362
rect 1846 348 1850 352
rect 1846 308 1850 312
rect 1814 268 1818 272
rect 1830 268 1834 272
rect 1790 258 1794 262
rect 1662 228 1666 232
rect 1782 228 1786 232
rect 1646 208 1650 212
rect 1742 198 1746 202
rect 1630 178 1634 182
rect 1622 148 1626 152
rect 1838 218 1842 222
rect 1862 278 1866 282
rect 1582 138 1586 142
rect 1614 138 1618 142
rect 1638 138 1642 142
rect 1726 138 1730 142
rect 1406 128 1410 132
rect 1438 128 1442 132
rect 1406 108 1410 112
rect 1278 88 1282 92
rect 1342 88 1346 92
rect 1366 88 1370 92
rect 1326 78 1330 82
rect 1302 68 1306 72
rect 1398 78 1402 82
rect 1382 68 1386 72
rect 1142 58 1146 62
rect 1270 58 1274 62
rect 1310 58 1314 62
rect 1142 48 1146 52
rect 862 38 866 42
rect 1126 38 1130 42
rect 1086 28 1090 32
rect 1342 28 1346 32
rect 1398 18 1402 22
rect 1430 18 1434 22
rect 1006 8 1010 12
rect 1198 8 1202 12
rect 1374 8 1378 12
rect 1418 3 1422 7
rect 1425 3 1429 7
rect 1566 128 1570 132
rect 1622 118 1626 122
rect 1598 108 1602 112
rect 1478 98 1482 102
rect 1622 98 1626 102
rect 1702 98 1706 102
rect 1726 98 1730 102
rect 1518 88 1522 92
rect 1502 78 1506 82
rect 1718 78 1722 82
rect 1942 588 1946 592
rect 1934 568 1938 572
rect 1918 558 1922 562
rect 1950 548 1954 552
rect 1958 548 1962 552
rect 1930 503 1934 507
rect 1937 503 1941 507
rect 1982 678 1986 682
rect 1974 658 1978 662
rect 1974 598 1978 602
rect 1998 738 2002 742
rect 2014 728 2018 732
rect 1998 718 2002 722
rect 2006 718 2010 722
rect 1998 598 2002 602
rect 1990 568 1994 572
rect 1982 558 1986 562
rect 1990 538 1994 542
rect 2366 1048 2370 1052
rect 2358 1008 2362 1012
rect 2366 998 2370 1002
rect 2358 958 2362 962
rect 2342 938 2346 942
rect 2366 938 2370 942
rect 2254 928 2258 932
rect 2350 928 2354 932
rect 2238 908 2242 912
rect 2310 898 2314 902
rect 2222 878 2226 882
rect 2166 868 2170 872
rect 2534 1098 2538 1102
rect 2542 1098 2546 1102
rect 2614 1178 2618 1182
rect 2622 1168 2626 1172
rect 2758 1258 2762 1262
rect 2710 1218 2714 1222
rect 2846 1328 2850 1332
rect 2854 1328 2858 1332
rect 2894 1328 2898 1332
rect 2806 1278 2810 1282
rect 2822 1278 2826 1282
rect 2870 1308 2874 1312
rect 2798 1268 2802 1272
rect 2838 1268 2842 1272
rect 2954 1503 2958 1507
rect 2961 1503 2965 1507
rect 3054 1518 3058 1522
rect 3038 1508 3042 1512
rect 3102 1478 3106 1482
rect 3086 1468 3090 1472
rect 3102 1468 3106 1472
rect 3190 1648 3194 1652
rect 3182 1638 3186 1642
rect 3142 1588 3146 1592
rect 3238 1808 3242 1812
rect 3254 1818 3258 1822
rect 3230 1748 3234 1752
rect 3246 1748 3250 1752
rect 3238 1738 3242 1742
rect 3222 1608 3226 1612
rect 3182 1578 3186 1582
rect 3142 1558 3146 1562
rect 3174 1558 3178 1562
rect 3134 1548 3138 1552
rect 3054 1458 3058 1462
rect 3126 1458 3130 1462
rect 3094 1448 3098 1452
rect 2998 1398 3002 1402
rect 3046 1398 3050 1402
rect 2926 1348 2930 1352
rect 2950 1348 2954 1352
rect 2934 1338 2938 1342
rect 2790 1258 2794 1262
rect 2870 1198 2874 1202
rect 2822 1168 2826 1172
rect 2774 1158 2778 1162
rect 2614 1148 2618 1152
rect 2630 1148 2634 1152
rect 2814 1148 2818 1152
rect 2574 1128 2578 1132
rect 2582 1128 2586 1132
rect 2614 1128 2618 1132
rect 2582 1108 2586 1112
rect 2462 1078 2466 1082
rect 2542 1078 2546 1082
rect 2478 1068 2482 1072
rect 2542 1068 2546 1072
rect 2478 1058 2482 1062
rect 2558 1058 2562 1062
rect 2382 1038 2386 1042
rect 2422 1038 2426 1042
rect 2430 1038 2434 1042
rect 2390 968 2394 972
rect 2486 1018 2490 1022
rect 2442 1003 2446 1007
rect 2449 1003 2453 1007
rect 2478 968 2482 972
rect 2518 998 2522 1002
rect 2502 958 2506 962
rect 2606 1088 2610 1092
rect 2638 1088 2642 1092
rect 2598 1078 2602 1082
rect 2966 1328 2970 1332
rect 2954 1303 2958 1307
rect 2961 1303 2965 1307
rect 2990 1278 2994 1282
rect 3022 1348 3026 1352
rect 3014 1338 3018 1342
rect 3038 1328 3042 1332
rect 3022 1308 3026 1312
rect 3030 1298 3034 1302
rect 3006 1268 3010 1272
rect 2998 1248 3002 1252
rect 3014 1218 3018 1222
rect 2990 1198 2994 1202
rect 3022 1198 3026 1202
rect 2910 1188 2914 1192
rect 2926 1188 2930 1192
rect 2894 1168 2898 1172
rect 2846 1158 2850 1162
rect 2854 1158 2858 1162
rect 2878 1158 2882 1162
rect 2894 1158 2898 1162
rect 2846 1148 2850 1152
rect 2870 1148 2874 1152
rect 2982 1178 2986 1182
rect 2934 1158 2938 1162
rect 2926 1148 2930 1152
rect 2934 1148 2938 1152
rect 2718 1118 2722 1122
rect 2734 1118 2738 1122
rect 2654 1078 2658 1082
rect 2678 1078 2682 1082
rect 2718 1078 2722 1082
rect 2670 1068 2674 1072
rect 2758 1068 2762 1072
rect 2622 1058 2626 1062
rect 2654 1058 2658 1062
rect 2774 1058 2778 1062
rect 2598 988 2602 992
rect 2542 978 2546 982
rect 2470 948 2474 952
rect 2510 948 2514 952
rect 2534 948 2538 952
rect 2406 938 2410 942
rect 2374 928 2378 932
rect 2398 928 2402 932
rect 2422 928 2426 932
rect 2382 918 2386 922
rect 2374 908 2378 912
rect 2622 968 2626 972
rect 2662 1048 2666 1052
rect 2686 1048 2690 1052
rect 2670 998 2674 1002
rect 2550 958 2554 962
rect 2630 958 2634 962
rect 2734 1008 2738 1012
rect 2758 978 2762 982
rect 2750 968 2754 972
rect 2790 968 2794 972
rect 2734 958 2738 962
rect 3006 1158 3010 1162
rect 2846 1118 2850 1122
rect 2862 1118 2866 1122
rect 2926 1118 2930 1122
rect 2950 1118 2954 1122
rect 2830 1098 2834 1102
rect 2894 1108 2898 1112
rect 2926 1098 2930 1102
rect 2954 1103 2958 1107
rect 2961 1103 2965 1107
rect 2862 1078 2866 1082
rect 2894 1078 2898 1082
rect 2918 1078 2922 1082
rect 2934 1078 2938 1082
rect 2958 1078 2962 1082
rect 2822 1068 2826 1072
rect 2870 1068 2874 1072
rect 2942 1068 2946 1072
rect 2854 988 2858 992
rect 2870 958 2874 962
rect 2894 988 2898 992
rect 3006 1128 3010 1132
rect 3014 1118 3018 1122
rect 2990 1098 2994 1102
rect 2934 1058 2938 1062
rect 2974 1058 2978 1062
rect 3006 1058 3010 1062
rect 2958 1048 2962 1052
rect 3006 1028 3010 1032
rect 2926 968 2930 972
rect 2894 958 2898 962
rect 2918 958 2922 962
rect 2630 948 2634 952
rect 2662 948 2666 952
rect 2766 948 2770 952
rect 2806 948 2810 952
rect 2814 948 2818 952
rect 2846 948 2850 952
rect 2470 938 2474 942
rect 2510 938 2514 942
rect 2622 938 2626 942
rect 2686 938 2690 942
rect 2734 938 2738 942
rect 2750 938 2754 942
rect 2446 928 2450 932
rect 2454 908 2458 912
rect 2430 878 2434 882
rect 2350 868 2354 872
rect 2398 868 2402 872
rect 2406 868 2410 872
rect 2422 868 2426 872
rect 2294 858 2298 862
rect 2302 858 2306 862
rect 2414 858 2418 862
rect 2438 858 2442 862
rect 2342 838 2346 842
rect 2366 838 2370 842
rect 2366 828 2370 832
rect 2310 818 2314 822
rect 2158 778 2162 782
rect 2206 778 2210 782
rect 2094 768 2098 772
rect 2302 778 2306 782
rect 2254 748 2258 752
rect 2294 748 2298 752
rect 2086 738 2090 742
rect 2158 738 2162 742
rect 2222 738 2226 742
rect 2078 728 2082 732
rect 2038 718 2042 722
rect 2174 728 2178 732
rect 2246 728 2250 732
rect 2086 698 2090 702
rect 2134 698 2138 702
rect 2182 698 2186 702
rect 2190 688 2194 692
rect 2094 678 2098 682
rect 2134 678 2138 682
rect 2022 608 2026 612
rect 2038 568 2042 572
rect 2022 548 2026 552
rect 2046 548 2050 552
rect 2054 538 2058 542
rect 2022 528 2026 532
rect 1950 498 1954 502
rect 2030 508 2034 512
rect 2006 488 2010 492
rect 2038 488 2042 492
rect 1950 468 1954 472
rect 1894 458 1898 462
rect 1894 448 1898 452
rect 1982 358 1986 362
rect 2006 438 2010 442
rect 2022 388 2026 392
rect 2006 358 2010 362
rect 1886 338 1890 342
rect 1934 338 1938 342
rect 1990 338 1994 342
rect 1998 328 2002 332
rect 1930 303 1934 307
rect 1937 303 1941 307
rect 1926 288 1930 292
rect 1878 278 1882 282
rect 1990 268 1994 272
rect 1870 258 1874 262
rect 2086 498 2090 502
rect 2118 558 2122 562
rect 2198 668 2202 672
rect 2230 668 2234 672
rect 2158 658 2162 662
rect 2222 658 2226 662
rect 2158 608 2162 612
rect 2142 588 2146 592
rect 2110 518 2114 522
rect 2134 518 2138 522
rect 2094 488 2098 492
rect 2150 558 2154 562
rect 2166 598 2170 602
rect 2158 548 2162 552
rect 2166 538 2170 542
rect 2158 478 2162 482
rect 2086 468 2090 472
rect 2078 448 2082 452
rect 2118 448 2122 452
rect 2126 448 2130 452
rect 2070 418 2074 422
rect 2094 418 2098 422
rect 2110 418 2114 422
rect 2102 408 2106 412
rect 2214 638 2218 642
rect 2230 638 2234 642
rect 2262 648 2266 652
rect 2254 638 2258 642
rect 2262 628 2266 632
rect 2246 578 2250 582
rect 2182 568 2186 572
rect 2222 568 2226 572
rect 2206 558 2210 562
rect 2214 548 2218 552
rect 2206 538 2210 542
rect 2182 528 2186 532
rect 2198 498 2202 502
rect 2174 468 2178 472
rect 2142 448 2146 452
rect 2150 438 2154 442
rect 2134 388 2138 392
rect 2166 348 2170 352
rect 2286 728 2290 732
rect 2278 718 2282 722
rect 2286 688 2290 692
rect 2302 678 2306 682
rect 2286 648 2290 652
rect 2294 648 2298 652
rect 2278 608 2282 612
rect 2278 568 2282 572
rect 2254 538 2258 542
rect 2294 538 2298 542
rect 2494 928 2498 932
rect 2510 918 2514 922
rect 2502 908 2506 912
rect 2486 888 2490 892
rect 2478 878 2482 882
rect 2494 878 2498 882
rect 2598 928 2602 932
rect 2534 918 2538 922
rect 2590 918 2594 922
rect 2566 898 2570 902
rect 2590 898 2594 902
rect 2646 918 2650 922
rect 2614 908 2618 912
rect 2614 898 2618 902
rect 2606 888 2610 892
rect 2518 878 2522 882
rect 2526 878 2530 882
rect 2582 878 2586 882
rect 2598 878 2602 882
rect 2574 868 2578 872
rect 2590 868 2594 872
rect 2518 858 2522 862
rect 2550 858 2554 862
rect 2462 848 2466 852
rect 2558 848 2562 852
rect 2494 838 2498 842
rect 2566 838 2570 842
rect 2574 838 2578 842
rect 2462 828 2466 832
rect 2414 818 2418 822
rect 2454 818 2458 822
rect 2326 758 2330 762
rect 2390 758 2394 762
rect 2318 698 2322 702
rect 2358 748 2362 752
rect 2398 748 2402 752
rect 2442 803 2446 807
rect 2449 803 2453 807
rect 2462 798 2466 802
rect 2430 778 2434 782
rect 2350 738 2354 742
rect 2390 738 2394 742
rect 2406 738 2410 742
rect 2318 688 2322 692
rect 2326 688 2330 692
rect 2366 708 2370 712
rect 2374 688 2378 692
rect 2350 678 2354 682
rect 2310 658 2314 662
rect 2334 658 2338 662
rect 2350 658 2354 662
rect 2342 648 2346 652
rect 2374 648 2378 652
rect 2310 638 2314 642
rect 2350 638 2354 642
rect 2262 518 2266 522
rect 2238 508 2242 512
rect 2254 488 2258 492
rect 2270 478 2274 482
rect 2286 398 2290 402
rect 2246 388 2250 392
rect 2350 618 2354 622
rect 2318 588 2322 592
rect 2350 568 2354 572
rect 2326 558 2330 562
rect 2318 538 2322 542
rect 2334 528 2338 532
rect 2422 708 2426 712
rect 2398 668 2402 672
rect 2382 598 2386 602
rect 2422 598 2426 602
rect 2406 578 2410 582
rect 2390 568 2394 572
rect 2398 558 2402 562
rect 2382 548 2386 552
rect 2342 518 2346 522
rect 2358 518 2362 522
rect 2422 498 2426 502
rect 2390 478 2394 482
rect 2406 468 2410 472
rect 2350 458 2354 462
rect 2326 448 2330 452
rect 2390 448 2394 452
rect 2254 358 2258 362
rect 2278 358 2282 362
rect 2310 358 2314 362
rect 2278 348 2282 352
rect 2294 348 2298 352
rect 2110 338 2114 342
rect 2038 328 2042 332
rect 2070 328 2074 332
rect 2126 308 2130 312
rect 2238 338 2242 342
rect 2078 298 2082 302
rect 2158 298 2162 302
rect 2206 298 2210 302
rect 2014 288 2018 292
rect 1886 228 1890 232
rect 1942 228 1946 232
rect 2022 268 2026 272
rect 2038 268 2042 272
rect 2070 268 2074 272
rect 2030 258 2034 262
rect 2014 218 2018 222
rect 1894 208 1898 212
rect 2022 178 2026 182
rect 1926 158 1930 162
rect 1950 158 1954 162
rect 1902 148 1906 152
rect 1958 148 1962 152
rect 1830 138 1834 142
rect 1894 138 1898 142
rect 1798 128 1802 132
rect 1814 118 1818 122
rect 1930 103 1934 107
rect 1937 103 1941 107
rect 1918 98 1922 102
rect 1790 88 1794 92
rect 1878 88 1882 92
rect 2046 228 2050 232
rect 2054 208 2058 212
rect 2038 158 2042 162
rect 2086 288 2090 292
rect 2094 288 2098 292
rect 2126 278 2130 282
rect 2166 288 2170 292
rect 2222 288 2226 292
rect 2142 268 2146 272
rect 2206 268 2210 272
rect 2086 218 2090 222
rect 2046 148 2050 152
rect 2062 148 2066 152
rect 2078 148 2082 152
rect 1998 138 2002 142
rect 2022 138 2026 142
rect 1974 128 1978 132
rect 2014 128 2018 132
rect 2006 118 2010 122
rect 1990 68 1994 72
rect 2014 68 2018 72
rect 2062 138 2066 142
rect 2086 138 2090 142
rect 2118 228 2122 232
rect 2134 218 2138 222
rect 2150 248 2154 252
rect 2262 318 2266 322
rect 2278 318 2282 322
rect 2278 298 2282 302
rect 2262 268 2266 272
rect 2318 348 2322 352
rect 2310 328 2314 332
rect 2366 428 2370 432
rect 2342 398 2346 402
rect 2334 368 2338 372
rect 2342 358 2346 362
rect 2334 338 2338 342
rect 2366 338 2370 342
rect 2382 338 2386 342
rect 2358 328 2362 332
rect 2374 328 2378 332
rect 2390 328 2394 332
rect 2382 298 2386 302
rect 2398 298 2402 302
rect 2366 288 2370 292
rect 2382 288 2386 292
rect 2310 278 2314 282
rect 2366 268 2370 272
rect 2230 248 2234 252
rect 2182 228 2186 232
rect 2174 198 2178 202
rect 2126 158 2130 162
rect 2110 148 2114 152
rect 2118 148 2122 152
rect 2142 148 2146 152
rect 2046 118 2050 122
rect 2094 118 2098 122
rect 2198 178 2202 182
rect 2190 158 2194 162
rect 2174 148 2178 152
rect 2182 148 2186 152
rect 2174 138 2178 142
rect 2158 98 2162 102
rect 2190 88 2194 92
rect 2062 78 2066 82
rect 2118 78 2122 82
rect 2150 78 2154 82
rect 2198 78 2202 82
rect 2166 68 2170 72
rect 2238 228 2242 232
rect 2230 188 2234 192
rect 2278 248 2282 252
rect 2446 758 2450 762
rect 2558 778 2562 782
rect 2478 758 2482 762
rect 2494 758 2498 762
rect 2438 748 2442 752
rect 2518 748 2522 752
rect 2502 728 2506 732
rect 2518 728 2522 732
rect 2470 708 2474 712
rect 2574 768 2578 772
rect 2582 748 2586 752
rect 2678 928 2682 932
rect 2710 918 2714 922
rect 2622 878 2626 882
rect 2670 878 2674 882
rect 2694 878 2698 882
rect 2830 928 2834 932
rect 2806 918 2810 922
rect 2806 908 2810 912
rect 2814 908 2818 912
rect 2830 908 2834 912
rect 2822 898 2826 902
rect 2822 878 2826 882
rect 2846 928 2850 932
rect 2870 928 2874 932
rect 2838 898 2842 902
rect 2878 888 2882 892
rect 2838 878 2842 882
rect 2662 868 2666 872
rect 2750 868 2754 872
rect 2782 868 2786 872
rect 2790 868 2794 872
rect 2622 858 2626 862
rect 2654 858 2658 862
rect 2766 858 2770 862
rect 2790 858 2794 862
rect 2630 828 2634 832
rect 2606 808 2610 812
rect 2606 768 2610 772
rect 2662 848 2666 852
rect 2638 808 2642 812
rect 2638 768 2642 772
rect 2582 738 2586 742
rect 2606 738 2610 742
rect 2614 738 2618 742
rect 2534 728 2538 732
rect 2558 728 2562 732
rect 2550 718 2554 722
rect 2486 698 2490 702
rect 2526 698 2530 702
rect 2590 708 2594 712
rect 2598 708 2602 712
rect 2614 708 2618 712
rect 2606 698 2610 702
rect 2502 678 2506 682
rect 2542 678 2546 682
rect 2478 608 2482 612
rect 2442 603 2446 607
rect 2449 603 2453 607
rect 2446 588 2450 592
rect 2806 848 2810 852
rect 2782 838 2786 842
rect 2774 828 2778 832
rect 2734 818 2738 822
rect 2742 818 2746 822
rect 2678 808 2682 812
rect 2686 808 2690 812
rect 2662 798 2666 802
rect 2678 798 2682 802
rect 2662 768 2666 772
rect 2670 748 2674 752
rect 2654 738 2658 742
rect 2654 728 2658 732
rect 2630 688 2634 692
rect 2646 688 2650 692
rect 2630 678 2634 682
rect 2614 668 2618 672
rect 2502 608 2506 612
rect 2486 598 2490 602
rect 2534 598 2538 602
rect 2606 658 2610 662
rect 2662 678 2666 682
rect 2670 678 2674 682
rect 2662 658 2666 662
rect 2910 928 2914 932
rect 2902 918 2906 922
rect 2926 898 2930 902
rect 3166 1548 3170 1552
rect 3214 1548 3218 1552
rect 3150 1528 3154 1532
rect 3182 1528 3186 1532
rect 3206 1528 3210 1532
rect 3158 1518 3162 1522
rect 3326 1858 3330 1862
rect 3310 1838 3314 1842
rect 3326 1838 3330 1842
rect 3278 1808 3282 1812
rect 3270 1778 3274 1782
rect 3278 1778 3282 1782
rect 3294 1758 3298 1762
rect 3526 1938 3530 1942
rect 3542 1928 3546 1932
rect 3574 1918 3578 1922
rect 3630 2038 3634 2042
rect 3654 2008 3658 2012
rect 3702 2268 3706 2272
rect 3710 2268 3714 2272
rect 3734 2268 3738 2272
rect 3782 2268 3786 2272
rect 3750 2258 3754 2262
rect 3782 2258 3786 2262
rect 3718 2238 3722 2242
rect 3726 2238 3730 2242
rect 3702 2218 3706 2222
rect 3678 2158 3682 2162
rect 3702 2158 3706 2162
rect 3702 2138 3706 2142
rect 3710 2098 3714 2102
rect 3678 2068 3682 2072
rect 3822 2258 3826 2262
rect 3814 2238 3818 2242
rect 3774 2228 3778 2232
rect 3822 2228 3826 2232
rect 3758 2208 3762 2212
rect 3734 2168 3738 2172
rect 3734 2158 3738 2162
rect 3758 2158 3762 2162
rect 3774 2158 3778 2162
rect 3806 2158 3810 2162
rect 3782 2148 3786 2152
rect 3862 2278 3866 2282
rect 3854 2268 3858 2272
rect 3838 2258 3842 2262
rect 3918 2298 3922 2302
rect 3910 2278 3914 2282
rect 3978 2303 3982 2307
rect 3985 2303 3989 2307
rect 3942 2298 3946 2302
rect 3982 2278 3986 2282
rect 3998 2278 4002 2282
rect 4014 2278 4018 2282
rect 4070 2318 4074 2322
rect 4086 2288 4090 2292
rect 4086 2278 4090 2282
rect 4166 2558 4170 2562
rect 4182 2668 4186 2672
rect 4150 2488 4154 2492
rect 4110 2458 4114 2462
rect 4134 2458 4138 2462
rect 4102 2368 4106 2372
rect 4118 2368 4122 2372
rect 4134 2358 4138 2362
rect 4118 2348 4122 2352
rect 4222 2738 4226 2742
rect 4238 2738 4242 2742
rect 4262 2728 4266 2732
rect 4270 2728 4274 2732
rect 4206 2718 4210 2722
rect 4254 2718 4258 2722
rect 4214 2678 4218 2682
rect 4262 2688 4266 2692
rect 4230 2648 4234 2652
rect 4222 2628 4226 2632
rect 4214 2568 4218 2572
rect 4190 2538 4194 2542
rect 4182 2488 4186 2492
rect 4158 2448 4162 2452
rect 4158 2418 4162 2422
rect 4174 2418 4178 2422
rect 4150 2368 4154 2372
rect 4318 2918 4322 2922
rect 4318 2898 4322 2902
rect 4310 2878 4314 2882
rect 4342 2948 4346 2952
rect 4350 2938 4354 2942
rect 4286 2818 4290 2822
rect 4302 2848 4306 2852
rect 4318 2848 4322 2852
rect 4310 2768 4314 2772
rect 4302 2758 4306 2762
rect 4358 2848 4362 2852
rect 4334 2748 4338 2752
rect 4310 2738 4314 2742
rect 4326 2738 4330 2742
rect 4334 2728 4338 2732
rect 4294 2718 4298 2722
rect 4326 2688 4330 2692
rect 4350 2708 4354 2712
rect 4382 2698 4386 2702
rect 4390 2698 4394 2702
rect 4390 2678 4394 2682
rect 4278 2668 4282 2672
rect 4286 2658 4290 2662
rect 4310 2658 4314 2662
rect 4342 2658 4346 2662
rect 4286 2648 4290 2652
rect 4342 2648 4346 2652
rect 4246 2578 4250 2582
rect 4270 2578 4274 2582
rect 4230 2548 4234 2552
rect 4350 2618 4354 2622
rect 4318 2548 4322 2552
rect 4366 2558 4370 2562
rect 4318 2528 4322 2532
rect 4358 2528 4362 2532
rect 4230 2478 4234 2482
rect 4374 2488 4378 2492
rect 4222 2468 4226 2472
rect 4302 2468 4306 2472
rect 4326 2468 4330 2472
rect 4358 2468 4362 2472
rect 4198 2388 4202 2392
rect 4182 2368 4186 2372
rect 4270 2458 4274 2462
rect 4294 2458 4298 2462
rect 4350 2458 4354 2462
rect 4294 2448 4298 2452
rect 4334 2448 4338 2452
rect 4238 2398 4242 2402
rect 4222 2358 4226 2362
rect 4230 2358 4234 2362
rect 4198 2348 4202 2352
rect 4150 2288 4154 2292
rect 4198 2338 4202 2342
rect 4222 2328 4226 2332
rect 4222 2318 4226 2322
rect 4214 2308 4218 2312
rect 4166 2278 4170 2282
rect 4174 2278 4178 2282
rect 4214 2278 4218 2282
rect 3942 2258 3946 2262
rect 3998 2258 4002 2262
rect 4022 2258 4026 2262
rect 4038 2258 4042 2262
rect 4054 2258 4058 2262
rect 3838 2248 3842 2252
rect 3934 2248 3938 2252
rect 3950 2248 3954 2252
rect 3846 2188 3850 2192
rect 3878 2238 3882 2242
rect 3886 2238 3890 2242
rect 3862 2198 3866 2202
rect 3854 2168 3858 2172
rect 3726 2138 3730 2142
rect 3750 2138 3754 2142
rect 3806 2138 3810 2142
rect 3838 2138 3842 2142
rect 3918 2218 3922 2222
rect 3910 2208 3914 2212
rect 3902 2198 3906 2202
rect 3958 2198 3962 2202
rect 4126 2248 4130 2252
rect 4142 2248 4146 2252
rect 4030 2238 4034 2242
rect 4062 2238 4066 2242
rect 3966 2168 3970 2172
rect 3950 2158 3954 2162
rect 3902 2148 3906 2152
rect 3758 2128 3762 2132
rect 3774 2128 3778 2132
rect 3822 2128 3826 2132
rect 3838 2128 3842 2132
rect 3854 2128 3858 2132
rect 3734 2118 3738 2122
rect 3718 2088 3722 2092
rect 3726 2088 3730 2092
rect 3806 2098 3810 2102
rect 3766 2078 3770 2082
rect 3790 2068 3794 2072
rect 3702 2058 3706 2062
rect 3718 2058 3722 2062
rect 3750 2058 3754 2062
rect 3702 2048 3706 2052
rect 3622 1988 3626 1992
rect 3622 1968 3626 1972
rect 3710 2038 3714 2042
rect 3758 2038 3762 2042
rect 3774 2048 3778 2052
rect 3830 2088 3834 2092
rect 3886 2128 3890 2132
rect 3878 2098 3882 2102
rect 3854 2078 3858 2082
rect 3846 2068 3850 2072
rect 4150 2188 4154 2192
rect 4134 2178 4138 2182
rect 4166 2168 4170 2172
rect 4062 2158 4066 2162
rect 4078 2158 4082 2162
rect 3926 2128 3930 2132
rect 3934 2088 3938 2092
rect 3918 2068 3922 2072
rect 3894 2058 3898 2062
rect 3814 2048 3818 2052
rect 3782 2028 3786 2032
rect 3910 2038 3914 2042
rect 3854 2018 3858 2022
rect 3758 1978 3762 1982
rect 3702 1958 3706 1962
rect 3590 1948 3594 1952
rect 3606 1948 3610 1952
rect 3622 1948 3626 1952
rect 3734 1948 3738 1952
rect 3670 1938 3674 1942
rect 3694 1938 3698 1942
rect 3718 1938 3722 1942
rect 3590 1928 3594 1932
rect 3630 1928 3634 1932
rect 3646 1928 3650 1932
rect 3510 1908 3514 1912
rect 3582 1908 3586 1912
rect 3446 1898 3450 1902
rect 3518 1898 3522 1902
rect 3430 1878 3434 1882
rect 3414 1868 3418 1872
rect 3542 1888 3546 1892
rect 3542 1878 3546 1882
rect 3558 1878 3562 1882
rect 3534 1868 3538 1872
rect 3550 1868 3554 1872
rect 3510 1858 3514 1862
rect 3374 1818 3378 1822
rect 3358 1808 3362 1812
rect 3382 1808 3386 1812
rect 3374 1778 3378 1782
rect 3366 1768 3370 1772
rect 3366 1758 3370 1762
rect 3278 1748 3282 1752
rect 3326 1748 3330 1752
rect 3350 1748 3354 1752
rect 3270 1738 3274 1742
rect 3294 1738 3298 1742
rect 3334 1738 3338 1742
rect 3310 1718 3314 1722
rect 3286 1708 3290 1712
rect 3374 1708 3378 1712
rect 3262 1698 3266 1702
rect 3310 1698 3314 1702
rect 3334 1698 3338 1702
rect 3254 1628 3258 1632
rect 3270 1608 3274 1612
rect 3262 1578 3266 1582
rect 3246 1558 3250 1562
rect 3254 1518 3258 1522
rect 3222 1498 3226 1502
rect 3238 1498 3242 1502
rect 3222 1478 3226 1482
rect 3166 1458 3170 1462
rect 3086 1408 3090 1412
rect 3070 1358 3074 1362
rect 3070 1288 3074 1292
rect 3054 1268 3058 1272
rect 3046 1258 3050 1262
rect 3070 1248 3074 1252
rect 3038 1198 3042 1202
rect 3038 1168 3042 1172
rect 3062 1158 3066 1162
rect 3230 1358 3234 1362
rect 3474 1803 3478 1807
rect 3481 1803 3485 1807
rect 3406 1768 3410 1772
rect 3430 1768 3434 1772
rect 3454 1758 3458 1762
rect 3462 1748 3466 1752
rect 3398 1738 3402 1742
rect 3430 1738 3434 1742
rect 3390 1718 3394 1722
rect 3406 1708 3410 1712
rect 3414 1698 3418 1702
rect 3414 1688 3418 1692
rect 3390 1678 3394 1682
rect 3406 1658 3410 1662
rect 3374 1628 3378 1632
rect 3294 1588 3298 1592
rect 3326 1588 3330 1592
rect 3286 1578 3290 1582
rect 3270 1558 3274 1562
rect 3310 1568 3314 1572
rect 3342 1568 3346 1572
rect 3294 1558 3298 1562
rect 3326 1558 3330 1562
rect 3366 1558 3370 1562
rect 3382 1608 3386 1612
rect 3382 1598 3386 1602
rect 3414 1588 3418 1592
rect 3406 1578 3410 1582
rect 3398 1568 3402 1572
rect 3374 1548 3378 1552
rect 3278 1528 3282 1532
rect 3334 1528 3338 1532
rect 3366 1528 3370 1532
rect 3374 1528 3378 1532
rect 3302 1518 3306 1522
rect 3350 1518 3354 1522
rect 3398 1558 3402 1562
rect 3414 1558 3418 1562
rect 3438 1718 3442 1722
rect 3446 1688 3450 1692
rect 3494 1678 3498 1682
rect 3438 1668 3442 1672
rect 3446 1658 3450 1662
rect 3462 1648 3466 1652
rect 3438 1628 3442 1632
rect 3446 1578 3450 1582
rect 3474 1603 3478 1607
rect 3481 1603 3485 1607
rect 3510 1738 3514 1742
rect 3510 1678 3514 1682
rect 3494 1588 3498 1592
rect 3470 1568 3474 1572
rect 3462 1558 3466 1562
rect 3622 1918 3626 1922
rect 3646 1898 3650 1902
rect 3598 1868 3602 1872
rect 3558 1858 3562 1862
rect 3606 1858 3610 1862
rect 3622 1858 3626 1862
rect 3678 1918 3682 1922
rect 3726 1918 3730 1922
rect 3702 1908 3706 1912
rect 3710 1888 3714 1892
rect 3742 1888 3746 1892
rect 3702 1878 3706 1882
rect 3742 1878 3746 1882
rect 3766 1878 3770 1882
rect 3598 1848 3602 1852
rect 3630 1848 3634 1852
rect 3534 1818 3538 1822
rect 3550 1798 3554 1802
rect 3598 1768 3602 1772
rect 3614 1758 3618 1762
rect 3590 1748 3594 1752
rect 3558 1738 3562 1742
rect 3550 1718 3554 1722
rect 3542 1708 3546 1712
rect 3582 1728 3586 1732
rect 3614 1728 3618 1732
rect 3566 1708 3570 1712
rect 3622 1708 3626 1712
rect 3646 1788 3650 1792
rect 3694 1858 3698 1862
rect 3678 1848 3682 1852
rect 3670 1838 3674 1842
rect 3846 2008 3850 2012
rect 3782 1938 3786 1942
rect 3918 1968 3922 1972
rect 3862 1948 3866 1952
rect 3894 1918 3898 1922
rect 3878 1908 3882 1912
rect 3806 1888 3810 1892
rect 3790 1878 3794 1882
rect 3862 1878 3866 1882
rect 3774 1868 3778 1872
rect 4054 2148 4058 2152
rect 4094 2148 4098 2152
rect 4102 2138 4106 2142
rect 4126 2138 4130 2142
rect 4286 2408 4290 2412
rect 4254 2398 4258 2402
rect 4318 2438 4322 2442
rect 4254 2348 4258 2352
rect 4310 2338 4314 2342
rect 4254 2308 4258 2312
rect 4286 2308 4290 2312
rect 4254 2288 4258 2292
rect 4262 2288 4266 2292
rect 4190 2268 4194 2272
rect 4198 2268 4202 2272
rect 4206 2268 4210 2272
rect 4246 2268 4250 2272
rect 4254 2268 4258 2272
rect 4182 2248 4186 2252
rect 4190 2158 4194 2162
rect 4158 2148 4162 2152
rect 4174 2148 4178 2152
rect 4198 2148 4202 2152
rect 4150 2138 4154 2142
rect 4062 2128 4066 2132
rect 4094 2128 4098 2132
rect 4134 2128 4138 2132
rect 4166 2128 4170 2132
rect 4126 2118 4130 2122
rect 4014 2108 4018 2112
rect 3978 2103 3982 2107
rect 3985 2103 3989 2107
rect 3998 2068 4002 2072
rect 3942 2058 3946 2062
rect 4078 2098 4082 2102
rect 4070 2078 4074 2082
rect 4022 2068 4026 2072
rect 4054 2068 4058 2072
rect 4014 2048 4018 2052
rect 4046 2038 4050 2042
rect 3950 2008 3954 2012
rect 4006 1958 4010 1962
rect 3958 1948 3962 1952
rect 4014 1948 4018 1952
rect 3934 1938 3938 1942
rect 3966 1938 3970 1942
rect 4078 1948 4082 1952
rect 4118 2078 4122 2082
rect 4102 2068 4106 2072
rect 4110 2058 4114 2062
rect 4118 2038 4122 2042
rect 4094 2028 4098 2032
rect 4094 1958 4098 1962
rect 4038 1938 4042 1942
rect 4070 1938 4074 1942
rect 4086 1938 4090 1942
rect 4014 1928 4018 1932
rect 4086 1928 4090 1932
rect 3902 1908 3906 1912
rect 3934 1898 3938 1902
rect 3758 1858 3762 1862
rect 3790 1858 3794 1862
rect 3822 1858 3826 1862
rect 3918 1858 3922 1862
rect 3734 1848 3738 1852
rect 3774 1848 3778 1852
rect 3978 1903 3982 1907
rect 3985 1903 3989 1907
rect 4006 1888 4010 1892
rect 3958 1878 3962 1882
rect 3942 1868 3946 1872
rect 3998 1868 4002 1872
rect 3942 1858 3946 1862
rect 3974 1858 3978 1862
rect 3990 1858 3994 1862
rect 3894 1848 3898 1852
rect 3774 1838 3778 1842
rect 3830 1838 3834 1842
rect 3718 1828 3722 1832
rect 3662 1818 3666 1822
rect 3742 1818 3746 1822
rect 3638 1768 3642 1772
rect 3750 1808 3754 1812
rect 3662 1778 3666 1782
rect 3726 1778 3730 1782
rect 3678 1758 3682 1762
rect 3734 1758 3738 1762
rect 3646 1708 3650 1712
rect 3606 1678 3610 1682
rect 3726 1748 3730 1752
rect 3758 1798 3762 1802
rect 3758 1778 3762 1782
rect 3766 1748 3770 1752
rect 3702 1738 3706 1742
rect 3774 1738 3778 1742
rect 3734 1718 3738 1722
rect 3702 1698 3706 1702
rect 3718 1698 3722 1702
rect 3686 1678 3690 1682
rect 3518 1668 3522 1672
rect 3574 1668 3578 1672
rect 3606 1668 3610 1672
rect 3622 1668 3626 1672
rect 3526 1658 3530 1662
rect 3518 1638 3522 1642
rect 3430 1548 3434 1552
rect 3462 1548 3466 1552
rect 3454 1528 3458 1532
rect 3430 1518 3434 1522
rect 3438 1518 3442 1522
rect 3302 1498 3306 1502
rect 3318 1488 3322 1492
rect 3302 1478 3306 1482
rect 3390 1498 3394 1502
rect 3422 1498 3426 1502
rect 3438 1488 3442 1492
rect 3334 1478 3338 1482
rect 3350 1478 3354 1482
rect 3382 1478 3386 1482
rect 3422 1478 3426 1482
rect 3294 1468 3298 1472
rect 3326 1468 3330 1472
rect 3342 1468 3346 1472
rect 3358 1468 3362 1472
rect 3374 1468 3378 1472
rect 3414 1468 3418 1472
rect 3278 1458 3282 1462
rect 3350 1448 3354 1452
rect 3414 1448 3418 1452
rect 3446 1448 3450 1452
rect 3382 1438 3386 1442
rect 3390 1438 3394 1442
rect 3406 1438 3410 1442
rect 3366 1398 3370 1402
rect 3278 1388 3282 1392
rect 3318 1368 3322 1372
rect 3430 1428 3434 1432
rect 3382 1368 3386 1372
rect 3342 1358 3346 1362
rect 3230 1348 3234 1352
rect 3262 1348 3266 1352
rect 3270 1348 3274 1352
rect 3398 1348 3402 1352
rect 3166 1328 3170 1332
rect 3150 1298 3154 1302
rect 3134 1288 3138 1292
rect 3150 1288 3154 1292
rect 3174 1288 3178 1292
rect 3126 1278 3130 1282
rect 3182 1268 3186 1272
rect 3254 1338 3258 1342
rect 3262 1298 3266 1302
rect 3238 1288 3242 1292
rect 3118 1248 3122 1252
rect 3158 1248 3162 1252
rect 3102 1218 3106 1222
rect 3094 1208 3098 1212
rect 3126 1208 3130 1212
rect 3214 1238 3218 1242
rect 3230 1238 3234 1242
rect 3174 1188 3178 1192
rect 3190 1178 3194 1182
rect 3150 1168 3154 1172
rect 3102 1158 3106 1162
rect 3134 1158 3138 1162
rect 3150 1158 3154 1162
rect 3166 1158 3170 1162
rect 3046 1148 3050 1152
rect 3078 1148 3082 1152
rect 3110 1148 3114 1152
rect 3078 1128 3082 1132
rect 3094 1128 3098 1132
rect 3118 1108 3122 1112
rect 3214 1188 3218 1192
rect 3222 1188 3226 1192
rect 3238 1188 3242 1192
rect 3254 1248 3258 1252
rect 3246 1178 3250 1182
rect 3262 1178 3266 1182
rect 3246 1158 3250 1162
rect 3198 1148 3202 1152
rect 3246 1148 3250 1152
rect 3190 1138 3194 1142
rect 3158 1128 3162 1132
rect 3134 1098 3138 1102
rect 3142 1098 3146 1102
rect 3110 1078 3114 1082
rect 3094 1068 3098 1072
rect 3182 1068 3186 1072
rect 3086 1008 3090 1012
rect 3110 1008 3114 1012
rect 3110 998 3114 1002
rect 3086 958 3090 962
rect 2942 918 2946 922
rect 3046 918 3050 922
rect 2954 903 2958 907
rect 2961 903 2965 907
rect 3054 898 3058 902
rect 2966 888 2970 892
rect 3046 888 3050 892
rect 2942 878 2946 882
rect 2854 868 2858 872
rect 2870 868 2874 872
rect 2894 868 2898 872
rect 2974 878 2978 882
rect 3078 878 3082 882
rect 2982 868 2986 872
rect 3006 868 3010 872
rect 2870 858 2874 862
rect 2894 848 2898 852
rect 2918 848 2922 852
rect 2950 848 2954 852
rect 2878 818 2882 822
rect 2814 798 2818 802
rect 2774 778 2778 782
rect 2774 748 2778 752
rect 2758 738 2762 742
rect 2894 808 2898 812
rect 2878 778 2882 782
rect 2846 768 2850 772
rect 2990 858 2994 862
rect 3102 908 3106 912
rect 3158 988 3162 992
rect 3118 968 3122 972
rect 3166 968 3170 972
rect 3126 948 3130 952
rect 3134 938 3138 942
rect 3142 938 3146 942
rect 3126 928 3130 932
rect 3110 888 3114 892
rect 3118 888 3122 892
rect 3142 888 3146 892
rect 3094 868 3098 872
rect 3134 868 3138 872
rect 3038 848 3042 852
rect 3070 848 3074 852
rect 3022 838 3026 842
rect 3054 828 3058 832
rect 3078 828 3082 832
rect 3038 798 3042 802
rect 3046 788 3050 792
rect 3046 778 3050 782
rect 2894 758 2898 762
rect 2966 758 2970 762
rect 2910 748 2914 752
rect 2926 748 2930 752
rect 2838 738 2842 742
rect 2862 738 2866 742
rect 2870 738 2874 742
rect 2710 728 2714 732
rect 2694 688 2698 692
rect 2718 718 2722 722
rect 2726 708 2730 712
rect 2790 678 2794 682
rect 2758 668 2762 672
rect 2798 668 2802 672
rect 2630 648 2634 652
rect 2574 588 2578 592
rect 2638 638 2642 642
rect 2590 558 2594 562
rect 2614 558 2618 562
rect 2686 578 2690 582
rect 2646 558 2650 562
rect 2670 558 2674 562
rect 2678 558 2682 562
rect 2590 548 2594 552
rect 2622 548 2626 552
rect 2478 538 2482 542
rect 2558 498 2562 502
rect 2518 488 2522 492
rect 2510 468 2514 472
rect 2534 468 2538 472
rect 2550 468 2554 472
rect 2462 458 2466 462
rect 2486 458 2490 462
rect 2462 408 2466 412
rect 2442 403 2446 407
rect 2449 403 2453 407
rect 2446 358 2450 362
rect 2414 338 2418 342
rect 2430 338 2434 342
rect 2406 288 2410 292
rect 2462 378 2466 382
rect 2502 448 2506 452
rect 2598 538 2602 542
rect 2614 538 2618 542
rect 2662 540 2666 544
rect 2750 658 2754 662
rect 2790 658 2794 662
rect 2758 648 2762 652
rect 2758 618 2762 622
rect 2750 598 2754 602
rect 2734 578 2738 582
rect 2718 558 2722 562
rect 2726 548 2730 552
rect 2742 548 2746 552
rect 2718 538 2722 542
rect 2582 458 2586 462
rect 2526 448 2530 452
rect 2534 448 2538 452
rect 2566 448 2570 452
rect 2590 448 2594 452
rect 2518 438 2522 442
rect 2582 398 2586 402
rect 2526 388 2530 392
rect 2478 368 2482 372
rect 2486 368 2490 372
rect 2510 368 2514 372
rect 2478 348 2482 352
rect 2502 348 2506 352
rect 2494 328 2498 332
rect 2486 308 2490 312
rect 2446 278 2450 282
rect 2494 278 2498 282
rect 2478 268 2482 272
rect 2558 378 2562 382
rect 2534 368 2538 372
rect 2542 348 2546 352
rect 2574 358 2578 362
rect 2566 348 2570 352
rect 2526 308 2530 312
rect 2534 298 2538 302
rect 2558 278 2562 282
rect 2518 268 2522 272
rect 2542 268 2546 272
rect 2398 258 2402 262
rect 2470 258 2474 262
rect 2510 258 2514 262
rect 2326 248 2330 252
rect 2350 248 2354 252
rect 2406 248 2410 252
rect 2406 238 2410 242
rect 2262 198 2266 202
rect 2286 198 2290 202
rect 2302 198 2306 202
rect 2254 168 2258 172
rect 2214 138 2218 142
rect 2230 138 2234 142
rect 2398 178 2402 182
rect 2286 148 2290 152
rect 2358 128 2362 132
rect 2342 118 2346 122
rect 2318 108 2322 112
rect 2350 108 2354 112
rect 2438 248 2442 252
rect 2478 248 2482 252
rect 2510 248 2514 252
rect 2462 218 2466 222
rect 2502 218 2506 222
rect 2526 218 2530 222
rect 2442 203 2446 207
rect 2449 203 2453 207
rect 2462 198 2466 202
rect 2494 198 2498 202
rect 2422 188 2426 192
rect 2414 138 2418 142
rect 2470 178 2474 182
rect 2502 178 2506 182
rect 2438 138 2442 142
rect 2462 138 2466 142
rect 2502 138 2506 142
rect 2382 78 2386 82
rect 2398 78 2402 82
rect 2486 128 2490 132
rect 2542 198 2546 202
rect 2534 178 2538 182
rect 2566 178 2570 182
rect 2558 148 2562 152
rect 2622 528 2626 532
rect 2630 518 2634 522
rect 2662 518 2666 522
rect 2606 448 2610 452
rect 2614 438 2618 442
rect 2622 358 2626 362
rect 2598 348 2602 352
rect 2702 518 2706 522
rect 2710 508 2714 512
rect 2678 498 2682 502
rect 2686 498 2690 502
rect 2702 488 2706 492
rect 2646 468 2650 472
rect 2734 468 2738 472
rect 2686 438 2690 442
rect 2638 408 2642 412
rect 2638 388 2642 392
rect 2654 378 2658 382
rect 2726 408 2730 412
rect 2702 388 2706 392
rect 2718 368 2722 372
rect 2686 358 2690 362
rect 2630 348 2634 352
rect 2662 348 2666 352
rect 2702 348 2706 352
rect 2606 338 2610 342
rect 2638 338 2642 342
rect 2702 338 2706 342
rect 2750 518 2754 522
rect 2774 578 2778 582
rect 2798 638 2802 642
rect 2790 608 2794 612
rect 2782 568 2786 572
rect 2822 708 2826 712
rect 2846 698 2850 702
rect 2854 678 2858 682
rect 2830 658 2834 662
rect 2822 648 2826 652
rect 2838 648 2842 652
rect 2822 558 2826 562
rect 2806 548 2810 552
rect 2782 538 2786 542
rect 2806 538 2810 542
rect 2854 588 2858 592
rect 2838 528 2842 532
rect 2822 518 2826 522
rect 2798 488 2802 492
rect 2798 478 2802 482
rect 2766 468 2770 472
rect 2766 458 2770 462
rect 2806 438 2810 442
rect 2766 398 2770 402
rect 2806 398 2810 402
rect 2734 348 2738 352
rect 2614 328 2618 332
rect 2678 328 2682 332
rect 2678 308 2682 312
rect 2622 298 2626 302
rect 2598 288 2602 292
rect 2590 268 2594 272
rect 2590 228 2594 232
rect 2582 198 2586 202
rect 2550 128 2554 132
rect 2566 128 2570 132
rect 2574 128 2578 132
rect 2534 118 2538 122
rect 2542 108 2546 112
rect 2486 78 2490 82
rect 2230 68 2234 72
rect 2254 68 2258 72
rect 2318 68 2322 72
rect 2590 178 2594 182
rect 2606 178 2610 182
rect 2686 288 2690 292
rect 2798 318 2802 322
rect 2742 288 2746 292
rect 2734 268 2738 272
rect 2798 308 2802 312
rect 2910 728 2914 732
rect 2926 728 2930 732
rect 2934 678 2938 682
rect 2886 668 2890 672
rect 2910 668 2914 672
rect 2982 748 2986 752
rect 3206 1128 3210 1132
rect 3198 1098 3202 1102
rect 3214 1078 3218 1082
rect 3230 1128 3234 1132
rect 3238 1118 3242 1122
rect 3246 1098 3250 1102
rect 3198 1058 3202 1062
rect 3222 1048 3226 1052
rect 3286 1338 3290 1342
rect 3294 1338 3298 1342
rect 3310 1338 3314 1342
rect 3342 1338 3346 1342
rect 3366 1338 3370 1342
rect 3334 1328 3338 1332
rect 3358 1328 3362 1332
rect 3294 1298 3298 1302
rect 3278 1268 3282 1272
rect 3310 1278 3314 1282
rect 3326 1278 3330 1282
rect 3358 1278 3362 1282
rect 3382 1278 3386 1282
rect 3390 1278 3394 1282
rect 3414 1298 3418 1302
rect 3278 1198 3282 1202
rect 3422 1288 3426 1292
rect 3350 1268 3354 1272
rect 3374 1268 3378 1272
rect 3406 1268 3410 1272
rect 3422 1268 3426 1272
rect 3318 1258 3322 1262
rect 3366 1258 3370 1262
rect 3310 1248 3314 1252
rect 3334 1248 3338 1252
rect 3350 1248 3354 1252
rect 3302 1228 3306 1232
rect 3358 1228 3362 1232
rect 3294 1188 3298 1192
rect 3286 1178 3290 1182
rect 3286 1168 3290 1172
rect 3334 1178 3338 1182
rect 3326 1158 3330 1162
rect 3382 1248 3386 1252
rect 3390 1238 3394 1242
rect 3398 1208 3402 1212
rect 3374 1198 3378 1202
rect 3406 1188 3410 1192
rect 3382 1168 3386 1172
rect 3278 1128 3282 1132
rect 3318 1128 3322 1132
rect 3350 1128 3354 1132
rect 3374 1128 3378 1132
rect 3286 1118 3290 1122
rect 3294 1118 3298 1122
rect 3262 1058 3266 1062
rect 3197 948 3201 952
rect 3198 918 3202 922
rect 3350 1108 3354 1112
rect 3342 1078 3346 1082
rect 3310 1068 3314 1072
rect 3334 1068 3338 1072
rect 3366 1068 3370 1072
rect 3342 1058 3346 1062
rect 3374 1058 3378 1062
rect 3414 1148 3418 1152
rect 3414 1128 3418 1132
rect 3398 1108 3402 1112
rect 3414 1068 3418 1072
rect 3454 1418 3458 1422
rect 3518 1528 3522 1532
rect 3526 1528 3530 1532
rect 3470 1518 3474 1522
rect 3494 1518 3498 1522
rect 3614 1658 3618 1662
rect 3550 1648 3554 1652
rect 3622 1648 3626 1652
rect 3606 1628 3610 1632
rect 3606 1608 3610 1612
rect 3646 1658 3650 1662
rect 3638 1598 3642 1602
rect 3646 1588 3650 1592
rect 3582 1578 3586 1582
rect 3926 1838 3930 1842
rect 3870 1818 3874 1822
rect 3894 1798 3898 1802
rect 3926 1798 3930 1802
rect 4022 1868 4026 1872
rect 3998 1848 4002 1852
rect 3950 1838 3954 1842
rect 4022 1798 4026 1802
rect 3950 1778 3954 1782
rect 3966 1778 3970 1782
rect 3942 1748 3946 1752
rect 3958 1748 3962 1752
rect 3838 1708 3842 1712
rect 3886 1708 3890 1712
rect 3934 1708 3938 1712
rect 3878 1698 3882 1702
rect 3830 1688 3834 1692
rect 3734 1678 3738 1682
rect 3758 1678 3762 1682
rect 3678 1658 3682 1662
rect 3734 1658 3738 1662
rect 3662 1648 3666 1652
rect 3694 1648 3698 1652
rect 3934 1658 3938 1662
rect 3958 1658 3962 1662
rect 3718 1648 3722 1652
rect 3846 1648 3850 1652
rect 3710 1638 3714 1642
rect 3942 1648 3946 1652
rect 3678 1608 3682 1612
rect 3678 1598 3682 1602
rect 3654 1568 3658 1572
rect 3662 1568 3666 1572
rect 3622 1558 3626 1562
rect 3638 1558 3642 1562
rect 3558 1548 3562 1552
rect 3590 1538 3594 1542
rect 3542 1528 3546 1532
rect 3574 1528 3578 1532
rect 3582 1528 3586 1532
rect 3598 1528 3602 1532
rect 3534 1518 3538 1522
rect 3558 1518 3562 1522
rect 3574 1508 3578 1512
rect 3534 1488 3538 1492
rect 3558 1478 3562 1482
rect 3670 1558 3674 1562
rect 3630 1538 3634 1542
rect 3654 1528 3658 1532
rect 3654 1508 3658 1512
rect 3838 1608 3842 1612
rect 3886 1608 3890 1612
rect 3814 1588 3818 1592
rect 3718 1578 3722 1582
rect 3790 1578 3794 1582
rect 3694 1568 3698 1572
rect 3686 1558 3690 1562
rect 3782 1558 3786 1562
rect 4070 1878 4074 1882
rect 4078 1878 4082 1882
rect 4150 2098 4154 2102
rect 4158 2068 4162 2072
rect 4142 2058 4146 2062
rect 4150 2038 4154 2042
rect 4134 2008 4138 2012
rect 4134 1968 4138 1972
rect 4198 2098 4202 2102
rect 4190 2088 4194 2092
rect 4174 2078 4178 2082
rect 4166 1978 4170 1982
rect 4214 2178 4218 2182
rect 4238 2258 4242 2262
rect 4230 2168 4234 2172
rect 4310 2298 4314 2302
rect 4390 2528 4394 2532
rect 4342 2438 4346 2442
rect 4382 2448 4386 2452
rect 4374 2368 4378 2372
rect 4342 2358 4346 2362
rect 4358 2358 4362 2362
rect 4382 2358 4386 2362
rect 4366 2348 4370 2352
rect 4326 2338 4330 2342
rect 4358 2318 4362 2322
rect 4350 2308 4354 2312
rect 4350 2298 4354 2302
rect 4318 2288 4322 2292
rect 4302 2278 4306 2282
rect 4294 2268 4298 2272
rect 4326 2278 4330 2282
rect 4262 2258 4266 2262
rect 4286 2258 4290 2262
rect 4262 2158 4266 2162
rect 4238 2148 4242 2152
rect 4222 2138 4226 2142
rect 4246 2118 4250 2122
rect 4278 2148 4282 2152
rect 4334 2268 4338 2272
rect 4374 2308 4378 2312
rect 4366 2278 4370 2282
rect 4350 2148 4354 2152
rect 4390 2228 4394 2232
rect 4382 2138 4386 2142
rect 4278 2128 4282 2132
rect 4270 2108 4274 2112
rect 4302 2118 4306 2122
rect 4294 2098 4298 2102
rect 4254 2078 4258 2082
rect 4262 2078 4266 2082
rect 4206 2068 4210 2072
rect 4246 2068 4250 2072
rect 4206 2048 4210 2052
rect 4382 2128 4386 2132
rect 4358 2098 4362 2102
rect 4326 2078 4330 2082
rect 4318 2068 4322 2072
rect 4334 2068 4338 2072
rect 4366 2068 4370 2072
rect 4358 2058 4362 2062
rect 4302 2048 4306 2052
rect 4270 2038 4274 2042
rect 4230 1998 4234 2002
rect 4214 1978 4218 1982
rect 4230 1968 4234 1972
rect 4302 2038 4306 2042
rect 4334 2038 4338 2042
rect 4294 1978 4298 1982
rect 4150 1958 4154 1962
rect 4270 1958 4274 1962
rect 4126 1948 4130 1952
rect 4142 1948 4146 1952
rect 4110 1938 4114 1942
rect 4166 1938 4170 1942
rect 4182 1938 4186 1942
rect 4198 1938 4202 1942
rect 4214 1938 4218 1942
rect 4158 1928 4162 1932
rect 4182 1928 4186 1932
rect 4222 1928 4226 1932
rect 4102 1908 4106 1912
rect 4150 1888 4154 1892
rect 4142 1868 4146 1872
rect 4078 1858 4082 1862
rect 4086 1858 4090 1862
rect 4110 1858 4114 1862
rect 4126 1858 4130 1862
rect 4062 1828 4066 1832
rect 4062 1818 4066 1822
rect 4046 1798 4050 1802
rect 4062 1798 4066 1802
rect 4038 1788 4042 1792
rect 4038 1768 4042 1772
rect 3974 1758 3978 1762
rect 3990 1758 3994 1762
rect 4006 1758 4010 1762
rect 4054 1758 4058 1762
rect 3998 1708 4002 1712
rect 3978 1703 3982 1707
rect 3985 1703 3989 1707
rect 4062 1708 4066 1712
rect 4086 1788 4090 1792
rect 4102 1788 4106 1792
rect 4102 1768 4106 1772
rect 4246 1898 4250 1902
rect 4230 1878 4234 1882
rect 4190 1868 4194 1872
rect 4150 1858 4154 1862
rect 4238 1858 4242 1862
rect 4174 1838 4178 1842
rect 4126 1798 4130 1802
rect 4126 1778 4130 1782
rect 4166 1828 4170 1832
rect 4278 1938 4282 1942
rect 4294 1948 4298 1952
rect 4302 1928 4306 1932
rect 4286 1918 4290 1922
rect 4302 1918 4306 1922
rect 4286 1908 4290 1912
rect 4278 1878 4282 1882
rect 4254 1858 4258 1862
rect 4198 1848 4202 1852
rect 4246 1848 4250 1852
rect 4198 1838 4202 1842
rect 4246 1838 4250 1842
rect 4158 1798 4162 1802
rect 4190 1788 4194 1792
rect 4206 1788 4210 1792
rect 4166 1778 4170 1782
rect 4158 1768 4162 1772
rect 4174 1768 4178 1772
rect 4118 1758 4122 1762
rect 4134 1758 4138 1762
rect 4142 1758 4146 1762
rect 4158 1758 4162 1762
rect 4182 1758 4186 1762
rect 4190 1758 4194 1762
rect 4094 1738 4098 1742
rect 4126 1748 4130 1752
rect 4134 1748 4138 1752
rect 4110 1718 4114 1722
rect 4102 1698 4106 1702
rect 4070 1678 4074 1682
rect 4078 1678 4082 1682
rect 4094 1668 4098 1672
rect 4006 1658 4010 1662
rect 4030 1658 4034 1662
rect 4054 1658 4058 1662
rect 4070 1658 4074 1662
rect 4142 1738 4146 1742
rect 4110 1658 4114 1662
rect 4134 1658 4138 1662
rect 4022 1648 4026 1652
rect 4078 1648 4082 1652
rect 4118 1648 4122 1652
rect 3942 1638 3946 1642
rect 3966 1638 3970 1642
rect 3950 1628 3954 1632
rect 3918 1578 3922 1582
rect 3862 1568 3866 1572
rect 4270 1828 4274 1832
rect 4342 1958 4346 1962
rect 4326 1938 4330 1942
rect 4366 1938 4370 1942
rect 4350 1928 4354 1932
rect 4358 1918 4362 1922
rect 4310 1908 4314 1912
rect 4310 1888 4314 1892
rect 4318 1868 4322 1872
rect 4334 1868 4338 1872
rect 4390 1928 4394 1932
rect 4366 1868 4370 1872
rect 4310 1858 4314 1862
rect 4358 1858 4362 1862
rect 4294 1828 4298 1832
rect 4278 1778 4282 1782
rect 4294 1778 4298 1782
rect 4326 1848 4330 1852
rect 4342 1848 4346 1852
rect 4214 1748 4218 1752
rect 4254 1748 4258 1752
rect 4190 1738 4194 1742
rect 4166 1728 4170 1732
rect 4190 1728 4194 1732
rect 4158 1718 4162 1722
rect 4174 1708 4178 1712
rect 4166 1668 4170 1672
rect 4150 1648 4154 1652
rect 4166 1648 4170 1652
rect 4182 1668 4186 1672
rect 4222 1728 4226 1732
rect 4214 1718 4218 1722
rect 4230 1718 4234 1722
rect 4230 1708 4234 1712
rect 4246 1708 4250 1712
rect 4222 1678 4226 1682
rect 4246 1688 4250 1692
rect 4198 1668 4202 1672
rect 4006 1638 4010 1642
rect 4062 1638 4066 1642
rect 4118 1638 4122 1642
rect 4142 1638 4146 1642
rect 4182 1638 4186 1642
rect 4014 1628 4018 1632
rect 4046 1628 4050 1632
rect 3998 1618 4002 1622
rect 4038 1578 4042 1582
rect 3822 1558 3826 1562
rect 3886 1558 3890 1562
rect 3926 1558 3930 1562
rect 3942 1558 3946 1562
rect 3990 1558 3994 1562
rect 4038 1558 4042 1562
rect 3686 1538 3690 1542
rect 3718 1538 3722 1542
rect 3734 1538 3738 1542
rect 3766 1538 3770 1542
rect 3798 1538 3802 1542
rect 3702 1528 3706 1532
rect 3742 1528 3746 1532
rect 3774 1528 3778 1532
rect 3718 1518 3722 1522
rect 3726 1518 3730 1522
rect 3718 1508 3722 1512
rect 3750 1508 3754 1512
rect 3606 1488 3610 1492
rect 3630 1488 3634 1492
rect 3606 1478 3610 1482
rect 3710 1478 3714 1482
rect 3470 1468 3474 1472
rect 3510 1468 3514 1472
rect 3566 1468 3570 1472
rect 3590 1468 3594 1472
rect 3622 1468 3626 1472
rect 3638 1468 3642 1472
rect 3694 1468 3698 1472
rect 3574 1458 3578 1462
rect 3550 1448 3554 1452
rect 3462 1408 3466 1412
rect 3438 1328 3442 1332
rect 3454 1298 3458 1302
rect 3474 1403 3478 1407
rect 3481 1403 3485 1407
rect 3550 1428 3554 1432
rect 3494 1398 3498 1402
rect 3526 1388 3530 1392
rect 3542 1368 3546 1372
rect 3734 1478 3738 1482
rect 3814 1518 3818 1522
rect 3766 1488 3770 1492
rect 3798 1488 3802 1492
rect 3782 1478 3786 1482
rect 3790 1478 3794 1482
rect 3670 1448 3674 1452
rect 3678 1448 3682 1452
rect 3582 1428 3586 1432
rect 3582 1418 3586 1422
rect 3598 1418 3602 1422
rect 3526 1328 3530 1332
rect 3478 1298 3482 1302
rect 3462 1278 3466 1282
rect 3438 1268 3442 1272
rect 3502 1288 3506 1292
rect 3534 1288 3538 1292
rect 3678 1438 3682 1442
rect 3734 1428 3738 1432
rect 3726 1408 3730 1412
rect 3702 1368 3706 1372
rect 3694 1358 3698 1362
rect 3614 1348 3618 1352
rect 3742 1408 3746 1412
rect 3750 1358 3754 1362
rect 3710 1348 3714 1352
rect 3606 1338 3610 1342
rect 3638 1338 3642 1342
rect 3654 1338 3658 1342
rect 3670 1338 3674 1342
rect 3654 1328 3658 1332
rect 3670 1328 3674 1332
rect 3694 1328 3698 1332
rect 3798 1468 3802 1472
rect 3790 1438 3794 1442
rect 3830 1478 3834 1482
rect 3902 1548 3906 1552
rect 3918 1538 3922 1542
rect 3934 1538 3938 1542
rect 3854 1518 3858 1522
rect 3998 1538 4002 1542
rect 3958 1528 3962 1532
rect 3942 1518 3946 1522
rect 3846 1508 3850 1512
rect 3902 1508 3906 1512
rect 3942 1488 3946 1492
rect 3978 1503 3982 1507
rect 3985 1503 3989 1507
rect 4006 1498 4010 1502
rect 4014 1498 4018 1502
rect 3838 1458 3842 1462
rect 3894 1458 3898 1462
rect 3822 1448 3826 1452
rect 3854 1448 3858 1452
rect 3806 1398 3810 1402
rect 3774 1358 3778 1362
rect 3806 1358 3810 1362
rect 3790 1348 3794 1352
rect 3734 1318 3738 1322
rect 3614 1288 3618 1292
rect 3686 1288 3690 1292
rect 3702 1288 3706 1292
rect 3726 1288 3730 1292
rect 3742 1288 3746 1292
rect 3614 1278 3618 1282
rect 3654 1278 3658 1282
rect 3694 1278 3698 1282
rect 3622 1268 3626 1272
rect 3670 1268 3674 1272
rect 3694 1258 3698 1262
rect 3510 1248 3514 1252
rect 3518 1248 3522 1252
rect 3494 1228 3498 1232
rect 3474 1203 3478 1207
rect 3481 1203 3485 1207
rect 3542 1248 3546 1252
rect 3582 1248 3586 1252
rect 3758 1288 3762 1292
rect 3782 1278 3786 1282
rect 3942 1438 3946 1442
rect 3854 1418 3858 1422
rect 3910 1408 3914 1412
rect 3902 1398 3906 1402
rect 3934 1398 3938 1402
rect 4054 1518 4058 1522
rect 4046 1508 4050 1512
rect 4022 1408 4026 1412
rect 3950 1378 3954 1382
rect 3958 1378 3962 1382
rect 4038 1378 4042 1382
rect 3838 1368 3842 1372
rect 3830 1358 3834 1362
rect 3870 1348 3874 1352
rect 3878 1338 3882 1342
rect 3806 1298 3810 1302
rect 3798 1288 3802 1292
rect 3814 1288 3818 1292
rect 3862 1288 3866 1292
rect 3878 1288 3882 1292
rect 3822 1278 3826 1282
rect 3750 1268 3754 1272
rect 3758 1268 3762 1272
rect 3790 1268 3794 1272
rect 3822 1268 3826 1272
rect 3974 1368 3978 1372
rect 4022 1358 4026 1362
rect 4118 1578 4122 1582
rect 4214 1618 4218 1622
rect 4222 1588 4226 1592
rect 4142 1568 4146 1572
rect 4198 1568 4202 1572
rect 4222 1568 4226 1572
rect 4086 1558 4090 1562
rect 4102 1558 4106 1562
rect 4102 1538 4106 1542
rect 4062 1508 4066 1512
rect 4070 1498 4074 1502
rect 4062 1478 4066 1482
rect 4054 1458 4058 1462
rect 4102 1468 4106 1472
rect 4118 1468 4122 1472
rect 4086 1448 4090 1452
rect 4110 1448 4114 1452
rect 4062 1438 4066 1442
rect 4078 1438 4082 1442
rect 4102 1438 4106 1442
rect 4086 1428 4090 1432
rect 4070 1378 4074 1382
rect 4062 1368 4066 1372
rect 4046 1358 4050 1362
rect 4078 1368 4082 1372
rect 3934 1348 3938 1352
rect 3950 1348 3954 1352
rect 3966 1348 3970 1352
rect 3990 1348 3994 1352
rect 4022 1348 4026 1352
rect 3918 1328 3922 1332
rect 3902 1308 3906 1312
rect 3894 1288 3898 1292
rect 3894 1268 3898 1272
rect 3830 1258 3834 1262
rect 3886 1258 3890 1262
rect 3606 1238 3610 1242
rect 3726 1238 3730 1242
rect 3526 1228 3530 1232
rect 3438 1178 3442 1182
rect 3454 1178 3458 1182
rect 3510 1178 3514 1182
rect 3590 1198 3594 1202
rect 3566 1188 3570 1192
rect 3526 1158 3530 1162
rect 3534 1158 3538 1162
rect 3438 1078 3442 1082
rect 3446 1068 3450 1072
rect 3446 1058 3450 1062
rect 3374 1048 3378 1052
rect 3286 1008 3290 1012
rect 3270 988 3274 992
rect 3350 1038 3354 1042
rect 3294 968 3298 972
rect 3238 958 3242 962
rect 3390 1008 3394 1012
rect 3294 948 3298 952
rect 3398 948 3402 952
rect 3326 928 3330 932
rect 3366 928 3370 932
rect 3262 908 3266 912
rect 3230 898 3234 902
rect 3182 888 3186 892
rect 3246 878 3250 882
rect 3222 868 3226 872
rect 3174 838 3178 842
rect 3174 828 3178 832
rect 3166 798 3170 802
rect 3134 768 3138 772
rect 3198 758 3202 762
rect 3150 748 3154 752
rect 3014 738 3018 742
rect 3038 738 3042 742
rect 2998 728 3002 732
rect 2990 718 2994 722
rect 3014 718 3018 722
rect 3070 718 3074 722
rect 3094 718 3098 722
rect 2954 703 2958 707
rect 2961 703 2965 707
rect 2966 688 2970 692
rect 2958 678 2962 682
rect 3022 688 3026 692
rect 3022 678 3026 682
rect 2974 668 2978 672
rect 3006 668 3010 672
rect 3134 708 3138 712
rect 3126 698 3130 702
rect 2998 658 3002 662
rect 3038 658 3042 662
rect 3062 658 3066 662
rect 2950 648 2954 652
rect 2982 648 2986 652
rect 3006 638 3010 642
rect 2910 628 2914 632
rect 2886 588 2890 592
rect 2878 578 2882 582
rect 3246 858 3250 862
rect 3230 848 3234 852
rect 3214 828 3218 832
rect 3222 798 3226 802
rect 3286 908 3290 912
rect 3278 898 3282 902
rect 3310 888 3314 892
rect 3262 848 3266 852
rect 3278 838 3282 842
rect 3246 788 3250 792
rect 3254 788 3258 792
rect 3294 768 3298 772
rect 3270 758 3274 762
rect 3318 808 3322 812
rect 3374 918 3378 922
rect 3382 908 3386 912
rect 3342 878 3346 882
rect 3374 878 3378 882
rect 3334 868 3338 872
rect 3422 938 3426 942
rect 3414 928 3418 932
rect 3406 908 3410 912
rect 3414 908 3418 912
rect 3342 858 3346 862
rect 3438 978 3442 982
rect 3494 1148 3498 1152
rect 3478 1138 3482 1142
rect 3462 1128 3466 1132
rect 3462 1108 3466 1112
rect 3470 1078 3474 1082
rect 3470 1048 3474 1052
rect 3478 1048 3482 1052
rect 3518 1118 3522 1122
rect 3518 1088 3522 1092
rect 3510 1078 3514 1082
rect 3670 1198 3674 1202
rect 3654 1188 3658 1192
rect 3702 1178 3706 1182
rect 3910 1288 3914 1292
rect 3926 1288 3930 1292
rect 3942 1288 3946 1292
rect 3918 1278 3922 1282
rect 3846 1248 3850 1252
rect 3926 1238 3930 1242
rect 4006 1328 4010 1332
rect 4030 1328 4034 1332
rect 3978 1303 3982 1307
rect 3985 1303 3989 1307
rect 3998 1268 4002 1272
rect 4022 1268 4026 1272
rect 4014 1258 4018 1262
rect 4046 1258 4050 1262
rect 4022 1248 4026 1252
rect 4038 1248 4042 1252
rect 3950 1238 3954 1242
rect 3934 1228 3938 1232
rect 3950 1218 3954 1222
rect 3750 1198 3754 1202
rect 3822 1208 3826 1212
rect 3806 1178 3810 1182
rect 3766 1168 3770 1172
rect 3702 1158 3706 1162
rect 3726 1158 3730 1162
rect 3758 1158 3762 1162
rect 3606 1148 3610 1152
rect 3622 1148 3626 1152
rect 3678 1148 3682 1152
rect 3718 1148 3722 1152
rect 3750 1148 3754 1152
rect 3694 1128 3698 1132
rect 3718 1128 3722 1132
rect 3558 1108 3562 1112
rect 3622 1108 3626 1112
rect 3550 1098 3554 1102
rect 3654 1098 3658 1102
rect 3566 1078 3570 1082
rect 3582 1078 3586 1082
rect 3622 1078 3626 1082
rect 3710 1108 3714 1112
rect 3726 1108 3730 1112
rect 3702 1088 3706 1092
rect 3670 1078 3674 1082
rect 3694 1078 3698 1082
rect 3846 1158 3850 1162
rect 3862 1158 3866 1162
rect 3774 1148 3778 1152
rect 3798 1148 3802 1152
rect 3766 1138 3770 1142
rect 3822 1138 3826 1142
rect 3742 1098 3746 1102
rect 3766 1088 3770 1092
rect 3814 1128 3818 1132
rect 3838 1128 3842 1132
rect 3886 1128 3890 1132
rect 3886 1118 3890 1122
rect 3838 1088 3842 1092
rect 3790 1078 3794 1082
rect 3598 1068 3602 1072
rect 3630 1068 3634 1072
rect 3654 1068 3658 1072
rect 3686 1068 3690 1072
rect 3718 1068 3722 1072
rect 3734 1068 3738 1072
rect 3510 1058 3514 1062
rect 3542 1058 3546 1062
rect 3574 1058 3578 1062
rect 3646 1058 3650 1062
rect 3662 1058 3666 1062
rect 3678 1058 3682 1062
rect 3790 1058 3794 1062
rect 3502 1048 3506 1052
rect 3494 1028 3498 1032
rect 3474 1003 3478 1007
rect 3481 1003 3485 1007
rect 3454 968 3458 972
rect 3598 1048 3602 1052
rect 3558 1038 3562 1042
rect 3662 1028 3666 1032
rect 3574 1008 3578 1012
rect 3534 988 3538 992
rect 3558 988 3562 992
rect 3518 968 3522 972
rect 3526 968 3530 972
rect 3510 958 3514 962
rect 3462 948 3466 952
rect 3478 948 3482 952
rect 3454 938 3458 942
rect 3462 928 3466 932
rect 3518 928 3522 932
rect 3446 918 3450 922
rect 3438 888 3442 892
rect 3422 878 3426 882
rect 3430 878 3434 882
rect 3430 868 3434 872
rect 3614 978 3618 982
rect 3598 958 3602 962
rect 3542 938 3546 942
rect 3550 928 3554 932
rect 3534 888 3538 892
rect 3462 868 3466 872
rect 3478 868 3482 872
rect 3366 858 3370 862
rect 3390 858 3394 862
rect 3398 858 3402 862
rect 3358 838 3362 842
rect 3422 828 3426 832
rect 3350 778 3354 782
rect 3286 748 3290 752
rect 3310 748 3314 752
rect 3510 858 3514 862
rect 3518 848 3522 852
rect 3470 838 3474 842
rect 3502 838 3506 842
rect 3474 803 3478 807
rect 3481 803 3485 807
rect 3494 798 3498 802
rect 3510 778 3514 782
rect 3454 758 3458 762
rect 3462 758 3466 762
rect 3494 758 3498 762
rect 3222 738 3226 742
rect 3278 738 3282 742
rect 3294 738 3298 742
rect 3310 728 3314 732
rect 3230 698 3234 702
rect 3110 628 3114 632
rect 3302 718 3306 722
rect 3238 688 3242 692
rect 3334 698 3338 702
rect 3422 718 3426 722
rect 3342 688 3346 692
rect 3358 688 3362 692
rect 3398 688 3402 692
rect 3406 688 3410 692
rect 3254 678 3258 682
rect 3270 678 3274 682
rect 3214 648 3218 652
rect 3254 648 3258 652
rect 3222 638 3226 642
rect 3062 588 3066 592
rect 3070 588 3074 592
rect 3086 588 3090 592
rect 3198 588 3202 592
rect 2926 548 2930 552
rect 2990 548 2994 552
rect 3174 578 3178 582
rect 3126 558 3130 562
rect 3166 558 3170 562
rect 3094 548 3098 552
rect 3118 548 3122 552
rect 3134 548 3138 552
rect 3150 548 3154 552
rect 2974 538 2978 542
rect 3118 538 3122 542
rect 3014 508 3018 512
rect 2954 503 2958 507
rect 2961 503 2965 507
rect 2934 498 2938 502
rect 2950 488 2954 492
rect 2878 478 2882 482
rect 2934 468 2938 472
rect 2974 358 2978 362
rect 3006 358 3010 362
rect 3062 478 3066 482
rect 3070 478 3074 482
rect 3094 478 3098 482
rect 3110 478 3114 482
rect 3038 468 3042 472
rect 3126 468 3130 472
rect 3190 558 3194 562
rect 3174 538 3178 542
rect 3230 608 3234 612
rect 3254 568 3258 572
rect 3230 558 3234 562
rect 3222 548 3226 552
rect 3214 538 3218 542
rect 3254 548 3258 552
rect 3238 538 3242 542
rect 3206 528 3210 532
rect 3230 518 3234 522
rect 3302 668 3306 672
rect 3334 668 3338 672
rect 3366 658 3370 662
rect 3390 658 3394 662
rect 3422 698 3426 702
rect 3382 648 3386 652
rect 3414 648 3418 652
rect 3526 768 3530 772
rect 3518 758 3522 762
rect 3534 728 3538 732
rect 3470 658 3474 662
rect 3494 658 3498 662
rect 3510 658 3514 662
rect 3454 638 3458 642
rect 3494 638 3498 642
rect 3286 588 3290 592
rect 3278 558 3282 562
rect 3270 538 3274 542
rect 3246 508 3250 512
rect 3166 478 3170 482
rect 3206 478 3210 482
rect 3166 468 3170 472
rect 3214 468 3218 472
rect 3230 468 3234 472
rect 3046 458 3050 462
rect 3078 458 3082 462
rect 3142 458 3146 462
rect 3158 458 3162 462
rect 3030 448 3034 452
rect 3094 448 3098 452
rect 3046 418 3050 422
rect 3062 358 3066 362
rect 2974 348 2978 352
rect 2998 348 3002 352
rect 2814 298 2818 302
rect 2846 298 2850 302
rect 2806 288 2810 292
rect 2806 278 2810 282
rect 2790 268 2794 272
rect 2750 258 2754 262
rect 2774 258 2778 262
rect 2702 248 2706 252
rect 2750 208 2754 212
rect 2646 198 2650 202
rect 2718 198 2722 202
rect 2630 178 2634 182
rect 2662 178 2666 182
rect 2726 178 2730 182
rect 2718 168 2722 172
rect 2686 158 2690 162
rect 2646 138 2650 142
rect 2614 128 2618 132
rect 2590 118 2594 122
rect 2638 128 2642 132
rect 2678 118 2682 122
rect 2638 108 2642 112
rect 2622 88 2626 92
rect 2670 88 2674 92
rect 2590 78 2594 82
rect 2606 78 2610 82
rect 2630 78 2634 82
rect 2662 78 2666 82
rect 2614 68 2618 72
rect 2678 78 2682 82
rect 2702 148 2706 152
rect 2822 238 2826 242
rect 2742 138 2746 142
rect 2774 138 2778 142
rect 2702 98 2706 102
rect 2702 88 2706 92
rect 2694 68 2698 72
rect 1446 58 1450 62
rect 1566 58 1570 62
rect 1662 58 1666 62
rect 1774 58 1778 62
rect 1782 58 1786 62
rect 1830 58 1834 62
rect 1894 58 1898 62
rect 1998 58 2002 62
rect 2054 58 2058 62
rect 2222 58 2226 62
rect 2278 58 2282 62
rect 2310 58 2314 62
rect 2342 58 2346 62
rect 2366 58 2370 62
rect 2654 58 2658 62
rect 2678 58 2682 62
rect 1598 48 1602 52
rect 2014 48 2018 52
rect 2022 38 2026 42
rect 2038 38 2042 42
rect 2158 38 2162 42
rect 2166 28 2170 32
rect 2134 8 2138 12
rect 2150 8 2154 12
rect 2766 128 2770 132
rect 2790 98 2794 102
rect 2782 78 2786 82
rect 2710 68 2714 72
rect 2830 208 2834 212
rect 2958 338 2962 342
rect 2942 308 2946 312
rect 2954 303 2958 307
rect 2961 303 2965 307
rect 2934 298 2938 302
rect 2942 288 2946 292
rect 2958 288 2962 292
rect 2870 248 2874 252
rect 2854 218 2858 222
rect 2950 208 2954 212
rect 2838 198 2842 202
rect 2870 168 2874 172
rect 2990 208 2994 212
rect 3014 338 3018 342
rect 3046 338 3050 342
rect 3022 298 3026 302
rect 3054 298 3058 302
rect 3110 408 3114 412
rect 3086 388 3090 392
rect 3078 378 3082 382
rect 3102 378 3106 382
rect 3078 338 3082 342
rect 3078 298 3082 302
rect 3030 288 3034 292
rect 3070 288 3074 292
rect 3062 268 3066 272
rect 3054 258 3058 262
rect 3078 258 3082 262
rect 3182 458 3186 462
rect 3238 458 3242 462
rect 3374 608 3378 612
rect 3430 608 3434 612
rect 3474 603 3478 607
rect 3481 603 3485 607
rect 3350 598 3354 602
rect 3334 588 3338 592
rect 3438 588 3442 592
rect 3310 568 3314 572
rect 3334 558 3338 562
rect 3302 548 3306 552
rect 3470 558 3474 562
rect 3542 678 3546 682
rect 3558 758 3562 762
rect 3566 758 3570 762
rect 3582 948 3586 952
rect 3622 948 3626 952
rect 3654 948 3658 952
rect 3606 918 3610 922
rect 3622 918 3626 922
rect 3638 918 3642 922
rect 3646 908 3650 912
rect 3622 888 3626 892
rect 3582 848 3586 852
rect 3646 798 3650 802
rect 3582 778 3586 782
rect 3654 778 3658 782
rect 3590 768 3594 772
rect 3614 768 3618 772
rect 3638 748 3642 752
rect 3598 738 3602 742
rect 3630 738 3634 742
rect 3558 728 3562 732
rect 3590 728 3594 732
rect 3614 728 3618 732
rect 3590 688 3594 692
rect 3558 678 3562 682
rect 3550 658 3554 662
rect 3526 648 3530 652
rect 3542 648 3546 652
rect 3310 538 3314 542
rect 3310 528 3314 532
rect 3510 528 3514 532
rect 3422 518 3426 522
rect 3302 508 3306 512
rect 3302 468 3306 472
rect 3278 458 3282 462
rect 3190 448 3194 452
rect 3198 448 3202 452
rect 3254 418 3258 422
rect 3214 398 3218 402
rect 3190 388 3194 392
rect 3174 378 3178 382
rect 3270 358 3274 362
rect 3286 348 3290 352
rect 3118 298 3122 302
rect 3150 288 3154 292
rect 3142 278 3146 282
rect 3110 268 3114 272
rect 3158 268 3162 272
rect 3134 258 3138 262
rect 3094 248 3098 252
rect 3046 238 3050 242
rect 3062 238 3066 242
rect 2998 188 3002 192
rect 3110 218 3114 222
rect 3062 158 3066 162
rect 3134 248 3138 252
rect 3126 148 3130 152
rect 2910 138 2914 142
rect 2934 138 2938 142
rect 2958 138 2962 142
rect 3054 138 3058 142
rect 2854 128 2858 132
rect 2870 118 2874 122
rect 2886 78 2890 82
rect 3142 128 3146 132
rect 2954 103 2958 107
rect 2961 103 2965 107
rect 3078 88 3082 92
rect 3006 78 3010 82
rect 3094 78 3098 82
rect 2966 68 2970 72
rect 2990 68 2994 72
rect 3254 338 3258 342
rect 3278 338 3282 342
rect 3294 338 3298 342
rect 3238 318 3242 322
rect 3302 318 3306 322
rect 3254 288 3258 292
rect 3406 488 3410 492
rect 3422 488 3426 492
rect 3566 648 3570 652
rect 3558 628 3562 632
rect 3574 628 3578 632
rect 3550 608 3554 612
rect 3534 568 3538 572
rect 3630 678 3634 682
rect 3614 658 3618 662
rect 3566 588 3570 592
rect 3598 588 3602 592
rect 3590 578 3594 582
rect 3574 568 3578 572
rect 3558 528 3562 532
rect 3582 518 3586 522
rect 3574 508 3578 512
rect 3582 508 3586 512
rect 3558 488 3562 492
rect 3518 458 3522 462
rect 3334 378 3338 382
rect 3414 378 3418 382
rect 3374 358 3378 362
rect 3326 348 3330 352
rect 3366 348 3370 352
rect 3390 348 3394 352
rect 3342 338 3346 342
rect 3318 318 3322 322
rect 3334 308 3338 312
rect 3310 298 3314 302
rect 3390 318 3394 322
rect 3350 298 3354 302
rect 3302 278 3306 282
rect 3334 278 3338 282
rect 3318 268 3322 272
rect 3238 248 3242 252
rect 3238 228 3242 232
rect 3214 188 3218 192
rect 3198 178 3202 182
rect 3182 138 3186 142
rect 3174 118 3178 122
rect 3174 108 3178 112
rect 3214 88 3218 92
rect 3222 78 3226 82
rect 3342 258 3346 262
rect 3302 148 3306 152
rect 3382 298 3386 302
rect 3374 258 3378 262
rect 3366 248 3370 252
rect 3286 138 3290 142
rect 3358 138 3362 142
rect 3246 128 3250 132
rect 3590 468 3594 472
rect 3566 438 3570 442
rect 3474 403 3478 407
rect 3481 403 3485 407
rect 3534 398 3538 402
rect 3430 388 3434 392
rect 3470 348 3474 352
rect 3414 288 3418 292
rect 3438 288 3442 292
rect 3398 278 3402 282
rect 3406 278 3410 282
rect 3398 268 3402 272
rect 3390 148 3394 152
rect 3518 318 3522 322
rect 3486 308 3490 312
rect 3598 458 3602 462
rect 3662 768 3666 772
rect 3702 1048 3706 1052
rect 3702 1038 3706 1042
rect 3822 998 3826 1002
rect 3854 998 3858 1002
rect 3718 988 3722 992
rect 3734 988 3738 992
rect 3798 988 3802 992
rect 3782 958 3786 962
rect 3694 918 3698 922
rect 3686 758 3690 762
rect 3854 968 3858 972
rect 3870 968 3874 972
rect 3758 948 3762 952
rect 3774 948 3778 952
rect 3838 948 3842 952
rect 3734 938 3738 942
rect 3750 938 3754 942
rect 3814 938 3818 942
rect 3710 928 3714 932
rect 3710 918 3714 922
rect 3806 928 3810 932
rect 3814 928 3818 932
rect 3742 918 3746 922
rect 3758 918 3762 922
rect 3790 918 3794 922
rect 3742 898 3746 902
rect 3718 878 3722 882
rect 3726 878 3730 882
rect 3734 878 3738 882
rect 3742 868 3746 872
rect 3790 908 3794 912
rect 3798 888 3802 892
rect 3782 878 3786 882
rect 3846 898 3850 902
rect 3822 878 3826 882
rect 3862 878 3866 882
rect 3766 868 3770 872
rect 3806 868 3810 872
rect 3878 958 3882 962
rect 3782 858 3786 862
rect 3814 858 3818 862
rect 3830 858 3834 862
rect 4094 1358 4098 1362
rect 4094 1348 4098 1352
rect 4142 1558 4146 1562
rect 4142 1468 4146 1472
rect 4158 1528 4162 1532
rect 4206 1548 4210 1552
rect 4174 1538 4178 1542
rect 4182 1538 4186 1542
rect 4214 1538 4218 1542
rect 4166 1518 4170 1522
rect 4206 1488 4210 1492
rect 4158 1478 4162 1482
rect 4190 1468 4194 1472
rect 4166 1458 4170 1462
rect 4166 1448 4170 1452
rect 4150 1438 4154 1442
rect 4214 1478 4218 1482
rect 4254 1678 4258 1682
rect 4270 1678 4274 1682
rect 4246 1658 4250 1662
rect 4262 1648 4266 1652
rect 4270 1638 4274 1642
rect 4286 1658 4290 1662
rect 4294 1648 4298 1652
rect 4294 1628 4298 1632
rect 4262 1578 4266 1582
rect 4270 1578 4274 1582
rect 4246 1558 4250 1562
rect 4230 1548 4234 1552
rect 4270 1548 4274 1552
rect 4294 1548 4298 1552
rect 4246 1538 4250 1542
rect 4286 1518 4290 1522
rect 4238 1498 4242 1502
rect 4238 1468 4242 1472
rect 4198 1438 4202 1442
rect 4214 1438 4218 1442
rect 4182 1428 4186 1432
rect 4222 1428 4226 1432
rect 4222 1398 4226 1402
rect 4190 1388 4194 1392
rect 4134 1378 4138 1382
rect 4166 1378 4170 1382
rect 4126 1358 4130 1362
rect 4150 1368 4154 1372
rect 4150 1358 4154 1362
rect 4182 1368 4186 1372
rect 4214 1368 4218 1372
rect 4118 1348 4122 1352
rect 4110 1328 4114 1332
rect 4126 1328 4130 1332
rect 4190 1328 4194 1332
rect 4102 1298 4106 1302
rect 4118 1298 4122 1302
rect 4086 1278 4090 1282
rect 4110 1238 4114 1242
rect 4110 1218 4114 1222
rect 4030 1208 4034 1212
rect 4062 1208 4066 1212
rect 4078 1208 4082 1212
rect 4030 1188 4034 1192
rect 3998 1178 4002 1182
rect 3974 1168 3978 1172
rect 4022 1168 4026 1172
rect 4054 1168 4058 1172
rect 3902 1158 3906 1162
rect 3926 1148 3930 1152
rect 3926 1138 3930 1142
rect 3934 1138 3938 1142
rect 3958 1138 3962 1142
rect 3902 1078 3906 1082
rect 3942 1108 3946 1112
rect 3942 1068 3946 1072
rect 3990 1158 3994 1162
rect 4062 1158 4066 1162
rect 4030 1148 4034 1152
rect 4070 1148 4074 1152
rect 4086 1148 4090 1152
rect 4006 1138 4010 1142
rect 4038 1138 4042 1142
rect 4070 1128 4074 1132
rect 4094 1128 4098 1132
rect 4206 1338 4210 1342
rect 4214 1338 4218 1342
rect 4182 1308 4186 1312
rect 4134 1248 4138 1252
rect 4134 1228 4138 1232
rect 4174 1218 4178 1222
rect 4198 1278 4202 1282
rect 4214 1268 4218 1272
rect 4278 1468 4282 1472
rect 4286 1448 4290 1452
rect 4262 1418 4266 1422
rect 4230 1388 4234 1392
rect 4318 1698 4322 1702
rect 4318 1658 4322 1662
rect 4342 1768 4346 1772
rect 4382 1828 4386 1832
rect 4366 1748 4370 1752
rect 4350 1688 4354 1692
rect 4358 1688 4362 1692
rect 4310 1608 4314 1612
rect 4358 1658 4362 1662
rect 4342 1648 4346 1652
rect 4334 1638 4338 1642
rect 4342 1628 4346 1632
rect 4334 1608 4338 1612
rect 4326 1578 4330 1582
rect 4318 1568 4322 1572
rect 4350 1618 4354 1622
rect 4358 1618 4362 1622
rect 4310 1548 4314 1552
rect 4342 1528 4346 1532
rect 4310 1488 4314 1492
rect 4310 1468 4314 1472
rect 4286 1368 4290 1372
rect 4286 1358 4290 1362
rect 4318 1458 4322 1462
rect 4342 1438 4346 1442
rect 4326 1418 4330 1422
rect 4350 1418 4354 1422
rect 4334 1358 4338 1362
rect 4342 1348 4346 1352
rect 4302 1338 4306 1342
rect 4254 1318 4258 1322
rect 4262 1318 4266 1322
rect 4286 1318 4290 1322
rect 4238 1308 4242 1312
rect 4246 1308 4250 1312
rect 4262 1308 4266 1312
rect 4230 1268 4234 1272
rect 4254 1268 4258 1272
rect 4358 1338 4362 1342
rect 4318 1328 4322 1332
rect 4286 1278 4290 1282
rect 4334 1278 4338 1282
rect 4270 1268 4274 1272
rect 4246 1258 4250 1262
rect 4262 1258 4266 1262
rect 4238 1208 4242 1212
rect 4190 1198 4194 1202
rect 4198 1198 4202 1202
rect 4182 1188 4186 1192
rect 4182 1168 4186 1172
rect 4350 1268 4354 1272
rect 4334 1258 4338 1262
rect 4326 1248 4330 1252
rect 4390 1758 4394 1762
rect 4374 1678 4378 1682
rect 4374 1658 4378 1662
rect 4374 1448 4378 1452
rect 4374 1378 4378 1382
rect 4390 1308 4394 1312
rect 4374 1278 4378 1282
rect 4358 1258 4362 1262
rect 4342 1238 4346 1242
rect 4358 1238 4362 1242
rect 4350 1198 4354 1202
rect 4214 1188 4218 1192
rect 4238 1188 4242 1192
rect 4262 1178 4266 1182
rect 4302 1178 4306 1182
rect 4326 1178 4330 1182
rect 4214 1168 4218 1172
rect 4342 1168 4346 1172
rect 4382 1188 4386 1192
rect 4366 1178 4370 1182
rect 4390 1178 4394 1182
rect 4366 1168 4370 1172
rect 4110 1158 4114 1162
rect 4118 1158 4122 1162
rect 4214 1158 4218 1162
rect 4310 1158 4314 1162
rect 4126 1148 4130 1152
rect 4150 1148 4154 1152
rect 3978 1103 3982 1107
rect 3985 1103 3989 1107
rect 4166 1138 4170 1142
rect 4198 1138 4202 1142
rect 4190 1128 4194 1132
rect 4158 1118 4162 1122
rect 3982 1088 3986 1092
rect 4174 1088 4178 1092
rect 3974 1068 3978 1072
rect 3942 1058 3946 1062
rect 3966 1058 3970 1062
rect 3966 1048 3970 1052
rect 4134 1078 4138 1082
rect 4198 1098 4202 1102
rect 4206 1088 4210 1092
rect 4198 1078 4202 1082
rect 4102 1068 4106 1072
rect 4150 1068 4154 1072
rect 4166 1068 4170 1072
rect 4190 1068 4194 1072
rect 4094 1058 4098 1062
rect 4142 1058 4146 1062
rect 4158 1058 4162 1062
rect 4182 1058 4186 1062
rect 4270 1128 4274 1132
rect 4262 1108 4266 1112
rect 4254 1098 4258 1102
rect 4294 1098 4298 1102
rect 4334 1148 4338 1152
rect 4358 1148 4362 1152
rect 4326 1138 4330 1142
rect 4326 1128 4330 1132
rect 4302 1078 4306 1082
rect 4310 1068 4314 1072
rect 4270 1058 4274 1062
rect 4286 1058 4290 1062
rect 4014 1048 4018 1052
rect 4046 1048 4050 1052
rect 4078 1048 4082 1052
rect 3966 988 3970 992
rect 3926 968 3930 972
rect 3926 948 3930 952
rect 3918 938 3922 942
rect 3950 938 3954 942
rect 3910 928 3914 932
rect 3998 1038 4002 1042
rect 4030 1038 4034 1042
rect 4006 1028 4010 1032
rect 4062 1038 4066 1042
rect 4094 1038 4098 1042
rect 4134 1038 4138 1042
rect 4094 1028 4098 1032
rect 4070 1018 4074 1022
rect 4038 1008 4042 1012
rect 4022 978 4026 982
rect 3990 948 3994 952
rect 3998 938 4002 942
rect 4070 998 4074 1002
rect 4150 1028 4154 1032
rect 4238 1048 4242 1052
rect 4270 1048 4274 1052
rect 4094 968 4098 972
rect 4030 948 4034 952
rect 4006 928 4010 932
rect 4022 928 4026 932
rect 3942 918 3946 922
rect 3982 918 3986 922
rect 3998 918 4002 922
rect 3978 903 3982 907
rect 3985 903 3989 907
rect 3942 878 3946 882
rect 3934 868 3938 872
rect 3766 848 3770 852
rect 3870 848 3874 852
rect 3750 828 3754 832
rect 3710 768 3714 772
rect 3742 768 3746 772
rect 3862 828 3866 832
rect 3886 818 3890 822
rect 3902 858 3906 862
rect 3910 858 3914 862
rect 3894 798 3898 802
rect 3822 778 3826 782
rect 3854 778 3858 782
rect 3846 768 3850 772
rect 3870 768 3874 772
rect 3934 848 3938 852
rect 4006 888 4010 892
rect 3998 858 4002 862
rect 4022 878 4026 882
rect 4014 868 4018 872
rect 3958 848 3962 852
rect 3974 848 3978 852
rect 4014 848 4018 852
rect 3918 838 3922 842
rect 3926 798 3930 802
rect 4094 958 4098 962
rect 4062 948 4066 952
rect 4046 938 4050 942
rect 4054 938 4058 942
rect 4038 928 4042 932
rect 4070 908 4074 912
rect 4062 898 4066 902
rect 4030 868 4034 872
rect 4118 948 4122 952
rect 4094 938 4098 942
rect 4126 938 4130 942
rect 4086 928 4090 932
rect 4078 898 4082 902
rect 4078 868 4082 872
rect 4006 838 4010 842
rect 4038 838 4042 842
rect 3966 828 3970 832
rect 4038 828 4042 832
rect 4126 898 4130 902
rect 4094 878 4098 882
rect 4118 878 4122 882
rect 4118 868 4122 872
rect 4206 1018 4210 1022
rect 4238 1038 4242 1042
rect 4230 1028 4234 1032
rect 4222 1018 4226 1022
rect 4270 1028 4274 1032
rect 4238 968 4242 972
rect 4246 968 4250 972
rect 4166 948 4170 952
rect 4182 918 4186 922
rect 4182 908 4186 912
rect 4158 898 4162 902
rect 4206 958 4210 962
rect 4254 958 4258 962
rect 4230 948 4234 952
rect 4254 948 4258 952
rect 4222 938 4226 942
rect 4246 938 4250 942
rect 4198 928 4202 932
rect 4222 928 4226 932
rect 4198 918 4202 922
rect 4190 888 4194 892
rect 4166 878 4170 882
rect 4174 878 4178 882
rect 4134 868 4138 872
rect 4142 848 4146 852
rect 4134 838 4138 842
rect 4110 828 4114 832
rect 4062 798 4066 802
rect 3990 788 3994 792
rect 4022 788 4026 792
rect 3942 778 3946 782
rect 3926 768 3930 772
rect 3934 768 3938 772
rect 3958 768 3962 772
rect 3790 758 3794 762
rect 3830 758 3834 762
rect 3926 758 3930 762
rect 3750 748 3754 752
rect 3806 748 3810 752
rect 3822 748 3826 752
rect 3854 748 3858 752
rect 3918 748 3922 752
rect 3926 748 3930 752
rect 3950 748 3954 752
rect 3702 728 3706 732
rect 3694 698 3698 702
rect 3678 678 3682 682
rect 3686 668 3690 672
rect 3670 658 3674 662
rect 3646 638 3650 642
rect 3614 558 3618 562
rect 3614 528 3618 532
rect 3638 608 3642 612
rect 3686 618 3690 622
rect 3678 608 3682 612
rect 3654 578 3658 582
rect 3678 578 3682 582
rect 3646 548 3650 552
rect 3638 538 3642 542
rect 3646 528 3650 532
rect 3638 498 3642 502
rect 3646 488 3650 492
rect 3630 458 3634 462
rect 3670 458 3674 462
rect 3598 448 3602 452
rect 3606 448 3610 452
rect 3718 678 3722 682
rect 3742 738 3746 742
rect 3790 738 3794 742
rect 3854 738 3858 742
rect 3782 728 3786 732
rect 3798 728 3802 732
rect 3742 698 3746 702
rect 3766 698 3770 702
rect 3798 698 3802 702
rect 3846 698 3850 702
rect 3750 678 3754 682
rect 3886 728 3890 732
rect 3910 728 3914 732
rect 3862 678 3866 682
rect 3870 678 3874 682
rect 3774 668 3778 672
rect 3806 668 3810 672
rect 3838 668 3842 672
rect 3718 658 3722 662
rect 3750 658 3754 662
rect 3774 658 3778 662
rect 3798 658 3802 662
rect 3822 658 3826 662
rect 3750 648 3754 652
rect 3710 608 3714 612
rect 3718 588 3722 592
rect 3702 568 3706 572
rect 3718 558 3722 562
rect 3774 558 3778 562
rect 3790 558 3794 562
rect 3742 548 3746 552
rect 3846 648 3850 652
rect 3830 638 3834 642
rect 3806 618 3810 622
rect 3806 568 3810 572
rect 3750 538 3754 542
rect 3662 448 3666 452
rect 3646 438 3650 442
rect 3654 398 3658 402
rect 3630 378 3634 382
rect 3646 378 3650 382
rect 3638 358 3642 362
rect 3678 388 3682 392
rect 3822 528 3826 532
rect 3846 528 3850 532
rect 3702 478 3706 482
rect 3694 468 3698 472
rect 3670 378 3674 382
rect 3686 378 3690 382
rect 3606 348 3610 352
rect 3678 338 3682 342
rect 3646 328 3650 332
rect 3606 318 3610 322
rect 3678 318 3682 322
rect 3590 308 3594 312
rect 3502 298 3506 302
rect 3558 298 3562 302
rect 3582 298 3586 302
rect 3526 288 3530 292
rect 3494 278 3498 282
rect 3518 278 3522 282
rect 3582 288 3586 292
rect 3574 278 3578 282
rect 3566 268 3570 272
rect 3542 258 3546 262
rect 3558 258 3562 262
rect 3638 288 3642 292
rect 3662 288 3666 292
rect 3598 278 3602 282
rect 3606 278 3610 282
rect 3622 278 3626 282
rect 3646 278 3650 282
rect 3726 418 3730 422
rect 3710 388 3714 392
rect 3718 358 3722 362
rect 3798 508 3802 512
rect 3814 508 3818 512
rect 3790 488 3794 492
rect 3766 478 3770 482
rect 3742 468 3746 472
rect 3766 468 3770 472
rect 3782 468 3786 472
rect 3774 458 3778 462
rect 3814 458 3818 462
rect 3822 448 3826 452
rect 3774 418 3778 422
rect 3798 408 3802 412
rect 3814 368 3818 372
rect 3878 668 3882 672
rect 3862 658 3866 662
rect 3886 658 3890 662
rect 3894 648 3898 652
rect 3934 588 3938 592
rect 4006 768 4010 772
rect 3998 758 4002 762
rect 3990 748 3994 752
rect 3966 708 3970 712
rect 3978 703 3982 707
rect 3985 703 3989 707
rect 4030 768 4034 772
rect 4046 768 4050 772
rect 4166 848 4170 852
rect 4158 818 4162 822
rect 4102 768 4106 772
rect 4062 738 4066 742
rect 4030 728 4034 732
rect 4014 718 4018 722
rect 4014 688 4018 692
rect 4006 658 4010 662
rect 4022 668 4026 672
rect 4046 658 4050 662
rect 4054 658 4058 662
rect 4118 758 4122 762
rect 4110 748 4114 752
rect 4166 738 4170 742
rect 4094 728 4098 732
rect 4126 728 4130 732
rect 4086 668 4090 672
rect 4070 648 4074 652
rect 4158 708 4162 712
rect 4190 868 4194 872
rect 4206 858 4210 862
rect 4230 858 4234 862
rect 4238 848 4242 852
rect 4190 818 4194 822
rect 4230 818 4234 822
rect 4238 778 4242 782
rect 4230 768 4234 772
rect 4174 678 4178 682
rect 4102 668 4106 672
rect 4126 668 4130 672
rect 4142 668 4146 672
rect 4118 658 4122 662
rect 3966 638 3970 642
rect 3982 638 3986 642
rect 4006 638 4010 642
rect 4070 638 4074 642
rect 4078 638 4082 642
rect 4086 638 4090 642
rect 3974 628 3978 632
rect 4054 628 4058 632
rect 4062 628 4066 632
rect 4030 578 4034 582
rect 4038 578 4042 582
rect 4062 578 4066 582
rect 3910 568 3914 572
rect 3942 568 3946 572
rect 3958 568 3962 572
rect 3990 568 3994 572
rect 3878 558 3882 562
rect 3894 558 3898 562
rect 3918 558 3922 562
rect 3902 548 3906 552
rect 3886 538 3890 542
rect 3838 478 3842 482
rect 3854 478 3858 482
rect 3870 478 3874 482
rect 3910 478 3914 482
rect 3878 468 3882 472
rect 3894 468 3898 472
rect 3838 448 3842 452
rect 3854 398 3858 402
rect 3854 378 3858 382
rect 3838 368 3842 372
rect 3862 368 3866 372
rect 3878 368 3882 372
rect 3846 358 3850 362
rect 3726 338 3730 342
rect 3734 338 3738 342
rect 3742 338 3746 342
rect 3726 328 3730 332
rect 3702 318 3706 322
rect 3694 278 3698 282
rect 3614 258 3618 262
rect 3478 248 3482 252
rect 3502 248 3506 252
rect 3566 248 3570 252
rect 3598 248 3602 252
rect 3406 178 3410 182
rect 3414 148 3418 152
rect 3374 138 3378 142
rect 3422 138 3426 142
rect 3438 128 3442 132
rect 3366 98 3370 102
rect 3342 88 3346 92
rect 3254 78 3258 82
rect 3158 68 3162 72
rect 3198 68 3202 72
rect 3214 68 3218 72
rect 3238 68 3242 72
rect 2758 58 2762 62
rect 2782 58 2786 62
rect 2814 58 2818 62
rect 2942 58 2946 62
rect 3038 58 3042 62
rect 3166 58 3170 62
rect 3182 58 3186 62
rect 3238 58 3242 62
rect 3334 58 3338 62
rect 2294 28 2298 32
rect 2310 18 2314 22
rect 2622 48 2626 52
rect 2638 48 2642 52
rect 2670 48 2674 52
rect 2742 48 2746 52
rect 3190 38 3194 42
rect 3270 48 3274 52
rect 3430 108 3434 112
rect 3474 203 3478 207
rect 3481 203 3485 207
rect 3470 168 3474 172
rect 3542 218 3546 222
rect 3454 98 3458 102
rect 3446 78 3450 82
rect 3558 208 3562 212
rect 3734 298 3738 302
rect 3718 278 3722 282
rect 3838 348 3842 352
rect 3822 338 3826 342
rect 3790 328 3794 332
rect 3950 558 3954 562
rect 3942 478 3946 482
rect 3966 558 3970 562
rect 3934 458 3938 462
rect 3926 428 3930 432
rect 3982 548 3986 552
rect 3998 508 4002 512
rect 3978 503 3982 507
rect 3985 503 3989 507
rect 4030 548 4034 552
rect 4014 488 4018 492
rect 3998 468 4002 472
rect 3990 448 3994 452
rect 3950 438 3954 442
rect 3966 428 3970 432
rect 3942 368 3946 372
rect 4142 628 4146 632
rect 4134 618 4138 622
rect 4102 588 4106 592
rect 4094 578 4098 582
rect 4174 648 4178 652
rect 4166 638 4170 642
rect 4086 568 4090 572
rect 4102 568 4106 572
rect 4134 568 4138 572
rect 4158 568 4162 572
rect 4198 748 4202 752
rect 4190 718 4194 722
rect 4222 748 4226 752
rect 4214 718 4218 722
rect 4206 688 4210 692
rect 4198 668 4202 672
rect 4222 658 4226 662
rect 4206 618 4210 622
rect 4270 938 4274 942
rect 4270 928 4274 932
rect 4254 898 4258 902
rect 4254 878 4258 882
rect 4286 918 4290 922
rect 4278 908 4282 912
rect 4342 1098 4346 1102
rect 4358 1098 4362 1102
rect 4358 1088 4362 1092
rect 4342 1068 4346 1072
rect 4302 1048 4306 1052
rect 4326 928 4330 932
rect 4270 848 4274 852
rect 4278 848 4282 852
rect 4318 898 4322 902
rect 4318 878 4322 882
rect 4302 858 4306 862
rect 4310 858 4314 862
rect 4374 1078 4378 1082
rect 4358 938 4362 942
rect 4350 878 4354 882
rect 4326 848 4330 852
rect 4294 838 4298 842
rect 4342 838 4346 842
rect 4326 828 4330 832
rect 4334 828 4338 832
rect 4366 838 4370 842
rect 4286 818 4290 822
rect 4326 818 4330 822
rect 4358 818 4362 822
rect 4302 808 4306 812
rect 4278 778 4282 782
rect 4310 768 4314 772
rect 4334 758 4338 762
rect 4374 758 4378 762
rect 4254 748 4258 752
rect 4302 748 4306 752
rect 4294 738 4298 742
rect 4238 678 4242 682
rect 4230 568 4234 572
rect 4070 558 4074 562
rect 4102 558 4106 562
rect 4134 558 4138 562
rect 4166 558 4170 562
rect 4182 558 4186 562
rect 4190 558 4194 562
rect 4062 548 4066 552
rect 4078 548 4082 552
rect 4110 548 4114 552
rect 4142 548 4146 552
rect 4174 548 4178 552
rect 4190 548 4194 552
rect 4046 518 4050 522
rect 4046 498 4050 502
rect 4038 468 4042 472
rect 4030 438 4034 442
rect 4014 358 4018 362
rect 3982 348 3986 352
rect 3854 338 3858 342
rect 3870 338 3874 342
rect 3894 338 3898 342
rect 3902 338 3906 342
rect 3998 338 4002 342
rect 3774 318 3778 322
rect 3814 298 3818 302
rect 3766 288 3770 292
rect 3790 288 3794 292
rect 3806 288 3810 292
rect 3806 278 3810 282
rect 3678 258 3682 262
rect 3726 258 3730 262
rect 3758 258 3762 262
rect 3630 248 3634 252
rect 3638 218 3642 222
rect 3630 188 3634 192
rect 3654 188 3658 192
rect 3622 168 3626 172
rect 3614 148 3618 152
rect 3614 138 3618 142
rect 3558 118 3562 122
rect 3534 88 3538 92
rect 3550 68 3554 72
rect 3606 98 3610 102
rect 3574 88 3578 92
rect 3582 88 3586 92
rect 3606 88 3610 92
rect 3710 248 3714 252
rect 3742 248 3746 252
rect 3806 268 3810 272
rect 3886 318 3890 322
rect 3798 258 3802 262
rect 3726 228 3730 232
rect 3766 228 3770 232
rect 3702 218 3706 222
rect 3718 208 3722 212
rect 3750 208 3754 212
rect 3678 198 3682 202
rect 3670 158 3674 162
rect 3662 118 3666 122
rect 3638 78 3642 82
rect 3646 78 3650 82
rect 3614 68 3618 72
rect 3790 248 3794 252
rect 3774 188 3778 192
rect 3734 158 3738 162
rect 3734 128 3738 132
rect 3718 118 3722 122
rect 3702 98 3706 102
rect 3710 88 3714 92
rect 3926 328 3930 332
rect 3934 328 3938 332
rect 3918 298 3922 302
rect 3918 278 3922 282
rect 3934 278 3938 282
rect 3966 328 3970 332
rect 3966 308 3970 312
rect 3978 303 3982 307
rect 3985 303 3989 307
rect 3982 288 3986 292
rect 4062 478 4066 482
rect 4102 468 4106 472
rect 4206 528 4210 532
rect 4214 528 4218 532
rect 4206 518 4210 522
rect 4158 478 4162 482
rect 4182 478 4186 482
rect 4206 478 4210 482
rect 4174 468 4178 472
rect 4366 748 4370 752
rect 4390 748 4394 752
rect 4342 728 4346 732
rect 4334 668 4338 672
rect 4318 658 4322 662
rect 4262 648 4266 652
rect 4262 618 4266 622
rect 4246 578 4250 582
rect 4270 608 4274 612
rect 4270 598 4274 602
rect 4294 648 4298 652
rect 4382 678 4386 682
rect 4374 668 4378 672
rect 4350 658 4354 662
rect 4294 638 4298 642
rect 4310 638 4314 642
rect 4326 638 4330 642
rect 4342 638 4346 642
rect 4366 608 4370 612
rect 4278 568 4282 572
rect 4310 568 4314 572
rect 4374 568 4378 572
rect 4254 558 4258 562
rect 4326 558 4330 562
rect 4278 548 4282 552
rect 4238 518 4242 522
rect 4238 488 4242 492
rect 4246 468 4250 472
rect 4294 538 4298 542
rect 4318 548 4322 552
rect 4302 508 4306 512
rect 4270 488 4274 492
rect 4294 478 4298 482
rect 4286 468 4290 472
rect 4054 458 4058 462
rect 4094 458 4098 462
rect 4150 458 4154 462
rect 4182 458 4186 462
rect 4222 458 4226 462
rect 4254 458 4258 462
rect 4278 458 4282 462
rect 4054 448 4058 452
rect 4086 448 4090 452
rect 4126 448 4130 452
rect 4174 448 4178 452
rect 4110 438 4114 442
rect 4126 438 4130 442
rect 4142 438 4146 442
rect 4094 428 4098 432
rect 4070 398 4074 402
rect 4230 438 4234 442
rect 4214 428 4218 432
rect 4206 418 4210 422
rect 4262 398 4266 402
rect 4310 468 4314 472
rect 4350 548 4354 552
rect 4358 548 4362 552
rect 4342 528 4346 532
rect 4342 458 4346 462
rect 4310 448 4314 452
rect 4326 448 4330 452
rect 4342 448 4346 452
rect 4326 438 4330 442
rect 4294 428 4298 432
rect 4318 428 4322 432
rect 4342 418 4346 422
rect 4366 458 4370 462
rect 4270 378 4274 382
rect 4198 368 4202 372
rect 4230 368 4234 372
rect 4262 368 4266 372
rect 4294 368 4298 372
rect 4326 368 4330 372
rect 4358 368 4362 372
rect 4166 358 4170 362
rect 4198 358 4202 362
rect 4230 358 4234 362
rect 4278 358 4282 362
rect 4294 358 4298 362
rect 4102 348 4106 352
rect 4190 348 4194 352
rect 4222 348 4226 352
rect 4254 348 4258 352
rect 4302 348 4306 352
rect 4086 338 4090 342
rect 4102 278 4106 282
rect 3894 268 3898 272
rect 4006 268 4010 272
rect 4078 268 4082 272
rect 3870 258 3874 262
rect 3886 258 3890 262
rect 3910 258 3914 262
rect 3934 258 3938 262
rect 3998 258 4002 262
rect 4014 258 4018 262
rect 4046 258 4050 262
rect 3846 238 3850 242
rect 3950 248 3954 252
rect 3918 238 3922 242
rect 3830 228 3834 232
rect 3870 228 3874 232
rect 3902 228 3906 232
rect 3894 198 3898 202
rect 3814 178 3818 182
rect 3862 178 3866 182
rect 3894 178 3898 182
rect 3814 158 3818 162
rect 3838 158 3842 162
rect 3854 158 3858 162
rect 3846 148 3850 152
rect 3838 138 3842 142
rect 3878 158 3882 162
rect 3926 158 3930 162
rect 3934 158 3938 162
rect 3902 148 3906 152
rect 3926 148 3930 152
rect 3982 238 3986 242
rect 4038 238 4042 242
rect 3998 228 4002 232
rect 4030 218 4034 222
rect 4046 208 4050 212
rect 3966 178 3970 182
rect 4350 348 4354 352
rect 4350 328 4354 332
rect 4334 308 4338 312
rect 4374 438 4378 442
rect 4366 318 4370 322
rect 4366 308 4370 312
rect 4198 288 4202 292
rect 4270 288 4274 292
rect 4182 278 4186 282
rect 4262 278 4266 282
rect 4286 278 4290 282
rect 4078 248 4082 252
rect 4070 228 4074 232
rect 4110 228 4114 232
rect 4086 198 4090 202
rect 4062 168 4066 172
rect 4110 168 4114 172
rect 4038 158 4042 162
rect 3974 148 3978 152
rect 4006 148 4010 152
rect 3878 138 3882 142
rect 3918 138 3922 142
rect 3942 128 3946 132
rect 3950 128 3954 132
rect 3790 118 3794 122
rect 3838 118 3842 122
rect 3806 98 3810 102
rect 3902 98 3906 102
rect 3686 68 3690 72
rect 3718 68 3722 72
rect 3978 103 3982 107
rect 3985 103 3989 107
rect 3966 88 3970 92
rect 3822 78 3826 82
rect 3958 78 3962 82
rect 4038 78 4042 82
rect 3878 68 3882 72
rect 4214 208 4218 212
rect 4206 178 4210 182
rect 4190 138 4194 142
rect 4126 128 4130 132
rect 4086 108 4090 112
rect 4134 108 4138 112
rect 4174 108 4178 112
rect 4070 68 4074 72
rect 4102 68 4106 72
rect 4142 78 4146 82
rect 4150 78 4154 82
rect 4174 78 4178 82
rect 4166 68 4170 72
rect 4286 258 4290 262
rect 4334 258 4338 262
rect 4294 228 4298 232
rect 4270 178 4274 182
rect 4286 168 4290 172
rect 4262 158 4266 162
rect 4262 118 4266 122
rect 4334 178 4338 182
rect 4318 158 4322 162
rect 4326 158 4330 162
rect 4302 148 4306 152
rect 4310 128 4314 132
rect 4302 118 4306 122
rect 4198 88 4202 92
rect 4246 78 4250 82
rect 4278 68 4282 72
rect 3966 58 3970 62
rect 4118 58 4122 62
rect 4206 58 4210 62
rect 3614 48 3618 52
rect 3638 48 3642 52
rect 3694 48 3698 52
rect 4318 68 4322 72
rect 3230 28 3234 32
rect 3374 28 3378 32
rect 3654 38 3658 42
rect 3670 38 3674 42
rect 4158 48 4162 52
rect 4390 168 4394 172
rect 4366 158 4370 162
rect 4374 128 4378 132
rect 4350 108 4354 112
rect 4358 98 4362 102
rect 4334 58 4338 62
rect 4174 38 4178 42
rect 2398 8 2402 12
rect 2566 8 2570 12
rect 2638 8 2642 12
rect 2750 8 2754 12
rect 4054 8 4058 12
rect 4070 8 4074 12
rect 2442 3 2446 7
rect 2449 3 2453 7
rect 3474 3 3478 7
rect 3481 3 3485 7
<< metal3 >>
rect 896 3103 898 3107
rect 902 3103 905 3107
rect 910 3103 912 3107
rect 1928 3103 1930 3107
rect 1934 3103 1937 3107
rect 1942 3103 1944 3107
rect 2952 3103 2954 3107
rect 2958 3103 2961 3107
rect 2966 3103 2968 3107
rect 3976 3103 3978 3107
rect 3982 3103 3985 3107
rect 3990 3103 3992 3107
rect 1138 3098 1142 3101
rect 1162 3098 1174 3101
rect 1202 3098 1254 3101
rect 1258 3098 1270 3101
rect 1338 3098 1358 3101
rect 1698 3098 1702 3101
rect 1898 3098 1902 3101
rect 1914 3098 1918 3101
rect 2178 3098 2182 3101
rect 2490 3098 2502 3101
rect 2610 3098 2638 3101
rect 1470 3092 1473 3098
rect 2142 3092 2145 3098
rect 2406 3092 2409 3098
rect 646 3088 654 3091
rect 658 3088 678 3091
rect 690 3088 838 3091
rect 3618 3088 3646 3091
rect 3650 3088 3862 3091
rect 4266 3088 4318 3091
rect 442 3078 566 3081
rect 602 3078 622 3081
rect 634 3078 718 3081
rect 1894 3081 1897 3088
rect 2510 3081 2513 3088
rect 1894 3078 3054 3081
rect 3506 3078 3558 3081
rect 3562 3078 3590 3081
rect 3594 3078 3678 3081
rect 3754 3078 3766 3081
rect 3858 3078 3886 3081
rect 4094 3081 4097 3088
rect 4094 3078 4150 3081
rect 4154 3078 4182 3081
rect 4202 3078 4286 3081
rect 214 3072 217 3078
rect 234 3068 454 3071
rect 554 3068 558 3071
rect 618 3068 654 3071
rect 658 3068 790 3071
rect 798 3071 801 3078
rect 798 3068 878 3071
rect 1054 3071 1057 3078
rect 954 3068 1057 3071
rect 1546 3068 2406 3071
rect 2410 3068 2670 3071
rect 3746 3068 3790 3071
rect 3826 3068 3926 3071
rect 3978 3068 4038 3071
rect 4090 3068 4142 3071
rect 4170 3068 4198 3071
rect 4234 3068 4238 3071
rect 4250 3068 4254 3071
rect 4282 3068 4286 3071
rect 34 3058 78 3061
rect 82 3058 230 3061
rect 314 3058 318 3061
rect 570 3058 582 3061
rect 626 3058 694 3061
rect 714 3058 734 3061
rect 738 3058 814 3061
rect 818 3058 838 3061
rect 1178 3058 1286 3061
rect 1602 3058 1606 3061
rect 1674 3058 1838 3061
rect 1850 3058 1878 3061
rect 2090 3058 2126 3061
rect 2666 3058 2726 3061
rect 2906 3058 2950 3061
rect 2954 3058 3086 3061
rect 3090 3058 3118 3061
rect 3234 3058 3294 3061
rect 3522 3058 3566 3061
rect 3626 3058 3670 3061
rect 3694 3061 3697 3068
rect 3674 3058 3697 3061
rect 3706 3058 3758 3061
rect 3882 3058 3902 3061
rect 4002 3058 4006 3061
rect 4026 3058 4062 3061
rect 4106 3058 4110 3061
rect 4162 3058 4302 3061
rect 182 3048 214 3051
rect 218 3048 310 3051
rect 314 3048 382 3051
rect 714 3048 753 3051
rect 834 3048 854 3051
rect 858 3048 958 3051
rect 2606 3051 2609 3058
rect 1114 3048 1137 3051
rect 2606 3048 3366 3051
rect 3370 3048 3382 3051
rect 3554 3048 3614 3051
rect 3690 3048 3766 3051
rect 3770 3048 3782 3051
rect 3802 3048 3830 3051
rect 3938 3048 3950 3051
rect 3954 3048 3998 3051
rect 4042 3048 4158 3051
rect 4162 3048 4174 3051
rect 4266 3048 4270 3051
rect 4298 3048 4302 3051
rect 182 3042 185 3048
rect 334 3042 337 3048
rect 750 3042 753 3048
rect 1134 3042 1137 3048
rect 4030 3042 4033 3048
rect 730 3038 734 3041
rect 946 3038 982 3041
rect 1138 3038 1174 3041
rect 1274 3038 2062 3041
rect 3058 3038 3190 3041
rect 3498 3038 3526 3041
rect 3530 3038 3654 3041
rect 3674 3038 3702 3041
rect 3722 3038 3766 3041
rect 3778 3038 3822 3041
rect 3866 3038 3894 3041
rect 3898 3038 3942 3041
rect 4114 3038 4174 3041
rect 4186 3038 4310 3041
rect 4110 3032 4113 3038
rect 546 3028 630 3031
rect 706 3028 926 3031
rect 1042 3028 1566 3031
rect 2282 3028 2606 3031
rect 3106 3028 3558 3031
rect 3570 3028 3609 3031
rect 3674 3028 4102 3031
rect 4130 3028 4190 3031
rect 4194 3028 4246 3031
rect 3606 3022 3609 3028
rect 10 3018 102 3021
rect 106 3018 1534 3021
rect 1962 3018 2086 3021
rect 2090 3018 2318 3021
rect 2442 3018 2470 3021
rect 3002 3018 3198 3021
rect 3458 3018 3526 3021
rect 3658 3018 3886 3021
rect 3890 3018 3910 3021
rect 3914 3018 3958 3021
rect 3962 3018 4166 3021
rect 4242 3018 4262 3021
rect 4294 3021 4297 3028
rect 4294 3018 4366 3021
rect 2674 3008 2926 3011
rect 3506 3008 3518 3011
rect 3522 3008 3718 3011
rect 3818 3008 4054 3011
rect 4146 3008 4294 3011
rect 392 3003 394 3007
rect 398 3003 401 3007
rect 406 3003 408 3007
rect 1416 3003 1418 3007
rect 1422 3003 1425 3007
rect 1430 3003 1432 3007
rect 2174 3002 2177 3008
rect 2440 3003 2442 3007
rect 2446 3003 2449 3007
rect 2454 3003 2456 3007
rect 3472 3003 3474 3007
rect 3478 3003 3481 3007
rect 3486 3003 3488 3007
rect 138 2998 262 3001
rect 2754 2998 2814 3001
rect 3714 2998 3878 3001
rect 3906 2998 3958 3001
rect 4050 2998 4142 3001
rect 4146 2998 4238 3001
rect 4250 2998 4262 3001
rect 4306 2998 4342 3001
rect 354 2988 478 2991
rect 482 2988 1030 2991
rect 1034 2988 1150 2991
rect 1154 2988 1182 2991
rect 1402 2988 1638 2991
rect 1798 2991 1801 2998
rect 1786 2988 1801 2991
rect 2034 2988 2046 2991
rect 2050 2988 2078 2991
rect 2194 2988 2542 2991
rect 3274 2988 3502 2991
rect 3562 2988 3670 2991
rect 3722 2988 3822 2991
rect 3834 2988 4001 2991
rect 4098 2988 4102 2991
rect 4218 2988 4374 2991
rect 3998 2982 4001 2988
rect 594 2978 622 2981
rect 626 2978 822 2981
rect 1346 2978 1537 2981
rect 1562 2978 1790 2981
rect 2514 2978 2566 2981
rect 3586 2978 3694 2981
rect 3770 2978 3854 2981
rect 4058 2978 4110 2981
rect 4202 2978 4374 2981
rect 1534 2972 1537 2978
rect 690 2968 878 2971
rect 938 2968 974 2971
rect 1482 2968 1486 2971
rect 2050 2968 2270 2971
rect 2274 2968 2422 2971
rect 2570 2968 2766 2971
rect 2802 2968 2806 2971
rect 2902 2971 2905 2978
rect 2874 2968 2905 2971
rect 3566 2971 3569 2978
rect 3210 2968 3569 2971
rect 3762 2968 3798 2971
rect 4090 2968 4118 2971
rect 4122 2968 4134 2971
rect 4154 2968 4166 2971
rect 4186 2968 4262 2971
rect 4330 2968 4334 2971
rect 862 2958 870 2961
rect 874 2958 990 2961
rect 1178 2958 1238 2961
rect 1582 2961 1585 2968
rect 3742 2962 3745 2968
rect 1538 2958 1585 2961
rect 1818 2958 2254 2961
rect 2282 2958 2294 2961
rect 2730 2958 2862 2961
rect 2866 2958 2913 2961
rect 2978 2958 3294 2961
rect 3426 2958 3438 2961
rect 3450 2958 3478 2961
rect 3482 2958 3489 2961
rect 3498 2958 3614 2961
rect 3626 2958 3638 2961
rect 3786 2958 3894 2961
rect 3946 2958 3950 2961
rect 4038 2961 4041 2968
rect 3962 2958 4041 2961
rect 4138 2958 4150 2961
rect 4154 2958 4174 2961
rect 4338 2958 4342 2961
rect 354 2948 374 2951
rect 386 2948 430 2951
rect 610 2948 614 2951
rect 618 2948 625 2951
rect 658 2948 678 2951
rect 1010 2948 1406 2951
rect 1462 2948 1465 2958
rect 2910 2952 2913 2958
rect 1482 2948 1577 2951
rect 1674 2948 1678 2951
rect 2090 2948 2182 2951
rect 2346 2948 2398 2951
rect 2402 2948 2470 2951
rect 2482 2948 2598 2951
rect 2658 2948 2758 2951
rect 2874 2948 2878 2951
rect 2914 2948 2998 2951
rect 3122 2948 3142 2951
rect 3146 2948 3158 2951
rect 3162 2948 3190 2951
rect 3226 2948 3406 2951
rect 3410 2948 3430 2951
rect 3482 2948 3654 2951
rect 3658 2948 3710 2951
rect 3986 2948 4022 2951
rect 4094 2951 4097 2958
rect 4190 2952 4193 2958
rect 4094 2948 4118 2951
rect 4122 2948 4150 2951
rect 4154 2948 4158 2951
rect 4226 2948 4254 2951
rect 4314 2948 4318 2951
rect 4366 2951 4369 2958
rect 4346 2948 4369 2951
rect 1574 2942 1577 2948
rect 3070 2942 3073 2948
rect 178 2938 350 2941
rect 546 2938 670 2941
rect 818 2938 830 2941
rect 834 2938 998 2941
rect 1002 2938 1086 2941
rect 1278 2938 1414 2941
rect 1434 2938 1470 2941
rect 1490 2938 1534 2941
rect 1626 2938 1694 2941
rect 1698 2938 2038 2941
rect 2066 2938 3070 2941
rect 3170 2938 3342 2941
rect 3442 2938 4070 2941
rect 4074 2938 4102 2941
rect 4106 2938 4350 2941
rect 426 2928 438 2931
rect 578 2928 622 2931
rect 626 2928 646 2931
rect 766 2931 769 2938
rect 1278 2932 1281 2938
rect 706 2928 769 2931
rect 786 2928 942 2931
rect 954 2928 1046 2931
rect 1394 2928 1478 2931
rect 1498 2928 1542 2931
rect 1574 2931 1577 2938
rect 1606 2931 1609 2938
rect 1574 2928 1609 2931
rect 1642 2928 1750 2931
rect 1754 2928 1966 2931
rect 2306 2928 2494 2931
rect 2562 2928 2673 2931
rect 2762 2928 2798 2931
rect 2810 2928 2838 2931
rect 2906 2928 2910 2931
rect 3210 2928 3278 2931
rect 3386 2928 3390 2931
rect 3410 2928 3414 2931
rect 3594 2928 3678 2931
rect 3690 2928 3694 2931
rect 3706 2928 3734 2931
rect 3738 2928 3758 2931
rect 3762 2928 3766 2931
rect 3842 2928 3926 2931
rect 4018 2928 4046 2931
rect 4050 2928 4086 2931
rect 4154 2928 4198 2931
rect 4210 2928 4214 2931
rect 4234 2928 4254 2931
rect 2166 2922 2169 2928
rect 2670 2922 2673 2928
rect 418 2918 558 2921
rect 562 2918 654 2921
rect 666 2918 902 2921
rect 906 2918 958 2921
rect 1250 2918 1294 2921
rect 1426 2918 1438 2921
rect 1442 2918 1510 2921
rect 1514 2918 1558 2921
rect 1570 2918 1582 2921
rect 1586 2918 1878 2921
rect 2450 2918 2566 2921
rect 2746 2918 2750 2921
rect 2786 2918 2846 2921
rect 2850 2918 2886 2921
rect 2890 2918 2942 2921
rect 2946 2918 3102 2921
rect 3282 2918 3366 2921
rect 3394 2918 3502 2921
rect 3642 2918 3726 2921
rect 3930 2918 3990 2921
rect 3994 2918 4222 2921
rect 4226 2918 4238 2921
rect 4258 2918 4286 2921
rect 4290 2918 4318 2921
rect 2582 2912 2585 2918
rect 66 2908 110 2911
rect 650 2908 854 2911
rect 930 2908 950 2911
rect 978 2908 1078 2911
rect 1082 2908 1486 2911
rect 1602 2908 1654 2911
rect 1698 2908 1702 2911
rect 1834 2908 1894 2911
rect 2042 2908 2174 2911
rect 2322 2908 2414 2911
rect 3378 2908 3542 2911
rect 3546 2908 3550 2911
rect 3714 2908 3934 2911
rect 4034 2908 4062 2911
rect 4066 2908 4134 2911
rect 4186 2908 4230 2911
rect 896 2903 898 2907
rect 902 2903 905 2907
rect 910 2903 912 2907
rect 1928 2903 1930 2907
rect 1934 2903 1937 2907
rect 1942 2903 1944 2907
rect 2952 2903 2954 2907
rect 2958 2903 2961 2907
rect 2966 2903 2968 2907
rect 3976 2903 3978 2907
rect 3982 2903 3985 2907
rect 3990 2903 3992 2907
rect 266 2898 358 2901
rect 362 2898 382 2901
rect 522 2898 542 2901
rect 546 2898 566 2901
rect 674 2898 838 2901
rect 930 2898 1142 2901
rect 1274 2898 1358 2901
rect 1402 2898 1430 2901
rect 1842 2898 1886 2901
rect 2034 2898 2054 2901
rect 2162 2898 2326 2901
rect 2330 2898 2414 2901
rect 2426 2898 2510 2901
rect 2586 2898 2822 2901
rect 2834 2898 2902 2901
rect 3058 2898 3078 2901
rect 3114 2898 3190 2901
rect 3322 2898 3334 2901
rect 3354 2898 3502 2901
rect 3538 2898 3593 2901
rect 3602 2898 3630 2901
rect 4002 2898 4166 2901
rect 4178 2898 4294 2901
rect 4298 2898 4318 2901
rect 434 2888 646 2891
rect 650 2888 934 2891
rect 946 2888 1014 2891
rect 1418 2888 1454 2891
rect 1482 2888 1542 2891
rect 1546 2888 1638 2891
rect 1954 2888 2558 2891
rect 2566 2888 2633 2891
rect 2890 2888 3126 2891
rect 3130 2888 3478 2891
rect 3490 2888 3494 2891
rect 3530 2888 3561 2891
rect 3578 2888 3582 2891
rect 3590 2891 3593 2898
rect 3718 2892 3721 2898
rect 3590 2888 3710 2891
rect 3770 2888 3790 2891
rect 3794 2888 3886 2891
rect 3938 2888 3966 2891
rect 4034 2888 4038 2891
rect 4042 2888 4206 2891
rect 282 2878 342 2881
rect 566 2878 574 2881
rect 578 2878 598 2881
rect 922 2878 1038 2881
rect 1066 2878 1438 2881
rect 1442 2878 1494 2881
rect 1722 2878 1742 2881
rect 1794 2878 2286 2881
rect 2338 2878 2526 2881
rect 2566 2881 2569 2888
rect 2630 2882 2633 2888
rect 2554 2878 2569 2881
rect 2578 2878 2614 2881
rect 2818 2878 2894 2881
rect 3234 2878 3278 2881
rect 3518 2881 3521 2888
rect 3558 2882 3561 2888
rect 3506 2878 3521 2881
rect 3546 2878 3550 2881
rect 3578 2878 3598 2881
rect 3602 2878 3638 2881
rect 3730 2878 3982 2881
rect 4010 2878 4097 2881
rect 4250 2878 4278 2881
rect 4282 2878 4286 2881
rect 4290 2878 4310 2881
rect 102 2872 105 2878
rect 3094 2872 3097 2878
rect 4094 2872 4097 2878
rect 554 2868 590 2871
rect 626 2868 662 2871
rect 882 2868 966 2871
rect 970 2868 1073 2871
rect 1202 2868 1206 2871
rect 1370 2868 1750 2871
rect 1778 2868 1814 2871
rect 1850 2868 2310 2871
rect 2314 2868 2838 2871
rect 3102 2868 3273 2871
rect 242 2858 262 2861
rect 478 2861 481 2868
rect 1070 2862 1073 2868
rect 1254 2862 1257 2868
rect 478 2858 502 2861
rect 554 2858 558 2861
rect 586 2858 766 2861
rect 882 2858 894 2861
rect 970 2858 1054 2861
rect 1450 2858 1462 2861
rect 1466 2858 1558 2861
rect 1658 2858 1838 2861
rect 1890 2858 1934 2861
rect 2154 2858 2158 2861
rect 2530 2858 2598 2861
rect 2866 2858 2950 2861
rect 3102 2861 3105 2868
rect 3270 2862 3273 2868
rect 3498 2868 3702 2871
rect 3706 2868 3782 2871
rect 3786 2868 3862 2871
rect 3890 2868 3910 2871
rect 3922 2868 3942 2871
rect 3962 2868 4006 2871
rect 4034 2868 4062 2871
rect 4130 2868 4134 2871
rect 4194 2868 4214 2871
rect 4250 2868 4270 2871
rect 3350 2862 3353 2868
rect 3862 2862 3865 2868
rect 2986 2858 3105 2861
rect 3202 2858 3246 2861
rect 3498 2858 3521 2861
rect 3530 2858 3550 2861
rect 3578 2858 3598 2861
rect 3618 2858 3654 2861
rect 3778 2858 3806 2861
rect 3810 2858 3838 2861
rect 3898 2858 3926 2861
rect 3970 2858 4014 2861
rect 4058 2858 4086 2861
rect 4122 2858 4142 2861
rect 4146 2858 4198 2861
rect 3518 2852 3521 2858
rect 574 2848 633 2851
rect 882 2848 929 2851
rect 574 2842 577 2848
rect 630 2842 633 2848
rect 926 2842 929 2848
rect 982 2848 1022 2851
rect 1378 2848 1385 2851
rect 1466 2848 1470 2851
rect 1682 2848 1774 2851
rect 1850 2848 2294 2851
rect 2298 2848 2462 2851
rect 2538 2848 2638 2851
rect 2642 2848 2750 2851
rect 2762 2848 3142 2851
rect 3146 2848 3190 2851
rect 3194 2848 3214 2851
rect 3266 2848 3494 2851
rect 3522 2848 3614 2851
rect 3618 2848 3678 2851
rect 3802 2848 3814 2851
rect 3818 2848 3854 2851
rect 3858 2848 3913 2851
rect 3954 2848 3974 2851
rect 4214 2851 4217 2858
rect 4034 2848 4270 2851
rect 4282 2848 4302 2851
rect 4322 2848 4358 2851
rect 982 2842 985 2848
rect 98 2838 534 2841
rect 1130 2838 1350 2841
rect 1382 2841 1385 2848
rect 3910 2842 3913 2848
rect 1382 2838 1670 2841
rect 1674 2838 1790 2841
rect 1794 2838 2486 2841
rect 2490 2838 3254 2841
rect 3546 2838 3574 2841
rect 3594 2838 3670 2841
rect 3842 2838 3886 2841
rect 3946 2838 4046 2841
rect 218 2828 246 2831
rect 250 2828 302 2831
rect 1374 2831 1377 2838
rect 1202 2828 1377 2831
rect 1506 2828 1782 2831
rect 1866 2828 2070 2831
rect 2346 2828 2350 2831
rect 2498 2828 2934 2831
rect 2938 2828 3254 2831
rect 3258 2828 3550 2831
rect 3554 2828 3614 2831
rect 3618 2828 3630 2831
rect 3642 2828 3838 2831
rect 3858 2828 3878 2831
rect 3882 2828 3934 2831
rect 158 2821 161 2828
rect 158 2818 470 2821
rect 474 2818 606 2821
rect 730 2818 742 2821
rect 1274 2818 1750 2821
rect 1754 2818 1982 2821
rect 2362 2818 2382 2821
rect 2442 2818 2465 2821
rect 2594 2818 2606 2821
rect 3458 2818 3574 2821
rect 3594 2818 3654 2821
rect 3706 2818 3918 2821
rect 4082 2818 4182 2821
rect 4186 2818 4286 2821
rect 1998 2812 2001 2818
rect 2462 2812 2465 2818
rect 2670 2812 2673 2818
rect 3006 2812 3009 2818
rect 258 2808 350 2811
rect 442 2808 526 2811
rect 530 2808 870 2811
rect 1186 2808 1222 2811
rect 1250 2808 1326 2811
rect 1330 2808 1382 2811
rect 1442 2808 1486 2811
rect 1490 2808 1742 2811
rect 1882 2808 1902 2811
rect 3410 2808 3446 2811
rect 3498 2808 3646 2811
rect 3746 2808 3774 2811
rect 3818 2808 3918 2811
rect 4210 2808 4246 2811
rect 392 2803 394 2807
rect 398 2803 401 2807
rect 406 2803 408 2807
rect 1416 2803 1418 2807
rect 1422 2803 1425 2807
rect 1430 2803 1432 2807
rect 2440 2803 2442 2807
rect 2446 2803 2449 2807
rect 2454 2803 2456 2807
rect 3472 2803 3474 2807
rect 3478 2803 3481 2807
rect 3486 2803 3488 2807
rect 506 2798 534 2801
rect 538 2798 694 2801
rect 698 2798 806 2801
rect 1130 2798 1150 2801
rect 1154 2798 1270 2801
rect 1778 2798 2062 2801
rect 2238 2798 2342 2801
rect 2346 2798 2414 2801
rect 3002 2798 3014 2801
rect 3066 2798 3134 2801
rect 3178 2798 3377 2801
rect 3554 2798 4038 2801
rect 4178 2798 4222 2801
rect 4226 2798 4358 2801
rect 34 2788 198 2791
rect 330 2788 422 2791
rect 466 2788 526 2791
rect 538 2788 1150 2791
rect 1530 2788 1542 2791
rect 2238 2791 2241 2798
rect 1826 2788 2241 2791
rect 2250 2788 2254 2791
rect 2346 2788 2750 2791
rect 2754 2788 2910 2791
rect 2922 2788 3366 2791
rect 3374 2791 3377 2798
rect 3374 2788 3510 2791
rect 3570 2788 3630 2791
rect 3802 2788 4030 2791
rect 4034 2788 4126 2791
rect 4146 2788 4150 2791
rect 18 2778 70 2781
rect 74 2778 174 2781
rect 362 2778 550 2781
rect 686 2778 1390 2781
rect 1874 2778 1886 2781
rect 1922 2778 3166 2781
rect 3330 2778 3886 2781
rect 3890 2778 3910 2781
rect 3914 2778 4006 2781
rect 4010 2778 4190 2781
rect 4194 2778 4214 2781
rect 686 2772 689 2778
rect 346 2768 537 2771
rect 858 2768 862 2771
rect 874 2768 950 2771
rect 954 2768 990 2771
rect 994 2768 1014 2771
rect 1258 2768 1646 2771
rect 1890 2768 1910 2771
rect 2218 2768 2262 2771
rect 2482 2768 2566 2771
rect 2594 2768 2622 2771
rect 2626 2768 2662 2771
rect 2666 2768 2734 2771
rect 2738 2768 2750 2771
rect 2810 2768 2918 2771
rect 3018 2768 3102 2771
rect 3434 2768 3446 2771
rect 3474 2768 3478 2771
rect 3658 2768 3790 2771
rect 3882 2768 4110 2771
rect 4290 2768 4310 2771
rect 22 2761 25 2768
rect 86 2762 89 2768
rect 534 2762 537 2768
rect 2094 2762 2097 2768
rect 22 2758 38 2761
rect 106 2758 158 2761
rect 162 2758 214 2761
rect 218 2758 462 2761
rect 482 2758 526 2761
rect 634 2758 670 2761
rect 722 2758 726 2761
rect 730 2758 758 2761
rect 826 2758 838 2761
rect 842 2758 910 2761
rect 1354 2758 1686 2761
rect 1690 2758 1710 2761
rect 1714 2758 1990 2761
rect 2202 2758 2302 2761
rect 2466 2758 3566 2761
rect 3570 2758 3582 2761
rect 3586 2758 3662 2761
rect 3666 2758 3942 2761
rect 3946 2758 4134 2761
rect 4138 2758 4198 2761
rect 4298 2758 4302 2761
rect 34 2748 166 2751
rect 170 2748 270 2751
rect 274 2748 310 2751
rect 422 2748 502 2751
rect 538 2748 574 2751
rect 586 2748 638 2751
rect 642 2748 734 2751
rect 754 2748 758 2751
rect 802 2748 806 2751
rect 834 2748 854 2751
rect 858 2748 870 2751
rect 890 2748 894 2751
rect 922 2748 998 2751
rect 1018 2748 1022 2751
rect 1050 2748 1054 2751
rect 1210 2748 1278 2751
rect 1474 2748 1494 2751
rect 1674 2748 1694 2751
rect 1698 2748 1750 2751
rect 2090 2748 2094 2751
rect 2134 2751 2137 2758
rect 2114 2748 2121 2751
rect 2134 2748 2158 2751
rect 2442 2748 2502 2751
rect 2546 2748 2582 2751
rect 2602 2748 2662 2751
rect 2666 2748 2678 2751
rect 2698 2748 2745 2751
rect 34 2738 38 2741
rect 58 2738 86 2741
rect 146 2738 241 2741
rect 250 2738 286 2741
rect 422 2741 425 2748
rect 2118 2742 2121 2748
rect 2230 2742 2233 2748
rect 2742 2742 2745 2748
rect 2754 2748 2798 2751
rect 2826 2748 2830 2751
rect 2834 2748 2886 2751
rect 3090 2748 3126 2751
rect 3138 2748 3166 2751
rect 3226 2748 3246 2751
rect 3402 2748 3446 2751
rect 3450 2748 3518 2751
rect 3546 2748 3550 2751
rect 3746 2748 3750 2751
rect 3786 2748 3798 2751
rect 3810 2748 3846 2751
rect 3874 2748 3894 2751
rect 3898 2748 3982 2751
rect 4186 2748 4198 2751
rect 4238 2751 4241 2758
rect 4238 2748 4246 2751
rect 4250 2748 4270 2751
rect 4274 2748 4334 2751
rect 2750 2742 2753 2748
rect 322 2738 425 2741
rect 430 2738 510 2741
rect 530 2738 534 2741
rect 746 2738 862 2741
rect 866 2738 966 2741
rect 978 2738 1006 2741
rect 1266 2738 1270 2741
rect 1614 2738 1622 2741
rect 1802 2738 1817 2741
rect 82 2728 102 2731
rect 106 2728 182 2731
rect 238 2731 241 2738
rect 430 2732 433 2738
rect 574 2732 577 2738
rect 1166 2732 1169 2738
rect 1614 2732 1617 2738
rect 1814 2732 1817 2738
rect 2006 2738 2054 2741
rect 2122 2738 2222 2741
rect 2538 2738 2561 2741
rect 2570 2738 2574 2741
rect 2650 2738 2654 2741
rect 2690 2738 2718 2741
rect 2786 2738 2806 2741
rect 2838 2738 2878 2741
rect 2882 2738 2934 2741
rect 3114 2738 3134 2741
rect 3382 2741 3385 2748
rect 3258 2738 3385 2741
rect 3494 2738 3502 2741
rect 3570 2738 3582 2741
rect 3646 2741 3649 2748
rect 3782 2741 3785 2748
rect 4062 2742 4065 2748
rect 3646 2738 3785 2741
rect 3834 2738 3838 2741
rect 4074 2738 4118 2741
rect 4170 2738 4222 2741
rect 4242 2738 4246 2741
rect 4282 2738 4310 2741
rect 4330 2738 4334 2741
rect 2006 2732 2009 2738
rect 2318 2732 2321 2738
rect 238 2728 278 2731
rect 414 2728 422 2731
rect 522 2728 534 2731
rect 610 2728 694 2731
rect 722 2728 782 2731
rect 810 2728 830 2731
rect 858 2728 910 2731
rect 914 2728 982 2731
rect 1218 2728 1334 2731
rect 2058 2728 2102 2731
rect 2146 2728 2150 2731
rect 2162 2728 2166 2731
rect 2558 2731 2561 2738
rect 2558 2728 2566 2731
rect 2730 2728 2753 2731
rect 2762 2728 2774 2731
rect 2838 2731 2841 2738
rect 3094 2732 3097 2738
rect 2778 2728 2841 2731
rect 2946 2728 2958 2731
rect 2994 2728 3001 2731
rect 3238 2731 3241 2738
rect 3202 2728 3241 2731
rect 3406 2731 3409 2738
rect 3494 2732 3497 2738
rect 3250 2728 3409 2731
rect 3418 2728 3422 2731
rect 3590 2728 3646 2731
rect 3650 2728 3694 2731
rect 3722 2728 3726 2731
rect 3738 2728 3758 2731
rect 3842 2728 3846 2731
rect 3874 2728 3934 2731
rect 3938 2728 3958 2731
rect 3970 2728 3974 2731
rect 4042 2728 4110 2731
rect 4114 2728 4118 2731
rect 4138 2728 4262 2731
rect 4274 2728 4334 2731
rect 414 2722 417 2728
rect 566 2722 569 2728
rect 1022 2722 1025 2728
rect 2598 2722 2601 2728
rect 2750 2722 2753 2728
rect 122 2718 174 2721
rect 178 2718 222 2721
rect 226 2718 326 2721
rect 570 2718 774 2721
rect 810 2718 862 2721
rect 866 2718 870 2721
rect 890 2718 950 2721
rect 954 2718 990 2721
rect 1170 2718 1206 2721
rect 1618 2718 1798 2721
rect 1914 2718 2270 2721
rect 2426 2718 2598 2721
rect 2846 2721 2849 2728
rect 2998 2722 3001 2728
rect 3590 2722 3593 2728
rect 2794 2718 2849 2721
rect 2914 2718 2918 2721
rect 3362 2718 3398 2721
rect 3466 2718 3534 2721
rect 3658 2718 3662 2721
rect 3698 2718 3702 2721
rect 3762 2718 3854 2721
rect 3970 2718 3982 2721
rect 4082 2718 4086 2721
rect 4098 2718 4126 2721
rect 4130 2718 4137 2721
rect 4258 2718 4294 2721
rect 4298 2718 4310 2721
rect 4206 2712 4209 2718
rect 98 2708 198 2711
rect 210 2708 302 2711
rect 306 2708 414 2711
rect 562 2708 750 2711
rect 754 2708 854 2711
rect 1138 2708 1142 2711
rect 1186 2708 1254 2711
rect 1490 2708 1918 2711
rect 2234 2708 2398 2711
rect 2410 2708 2542 2711
rect 2586 2708 2702 2711
rect 2706 2708 2838 2711
rect 3122 2708 3254 2711
rect 3386 2708 3502 2711
rect 3506 2708 3526 2711
rect 3530 2708 3598 2711
rect 3610 2708 3902 2711
rect 4002 2708 4054 2711
rect 4058 2708 4174 2711
rect 4234 2708 4350 2711
rect 896 2703 898 2707
rect 902 2703 905 2707
rect 910 2703 912 2707
rect 1046 2702 1049 2708
rect 1928 2703 1930 2707
rect 1934 2703 1937 2707
rect 1942 2703 1944 2707
rect 2952 2703 2954 2707
rect 2958 2703 2961 2707
rect 2966 2703 2968 2707
rect 3976 2703 3978 2707
rect 3982 2703 3985 2707
rect 3990 2703 3992 2707
rect 66 2698 422 2701
rect 554 2698 566 2701
rect 682 2698 814 2701
rect 1154 2698 1206 2701
rect 1562 2698 1582 2701
rect 2362 2698 2526 2701
rect 2530 2698 2542 2701
rect 2626 2698 2630 2701
rect 2698 2698 2734 2701
rect 2738 2698 2830 2701
rect 2834 2698 2862 2701
rect 3002 2698 3046 2701
rect 3050 2698 3110 2701
rect 3586 2698 3678 2701
rect 3682 2698 3710 2701
rect 4002 2698 4182 2701
rect 4186 2698 4374 2701
rect 4382 2692 4385 2698
rect 4390 2692 4393 2698
rect 202 2688 230 2691
rect 234 2688 478 2691
rect 482 2688 846 2691
rect 858 2688 870 2691
rect 874 2688 878 2691
rect 890 2688 894 2691
rect 1266 2688 1430 2691
rect 1634 2688 1686 2691
rect 1926 2688 2110 2691
rect 2114 2688 2222 2691
rect 2322 2688 2401 2691
rect 2426 2688 2582 2691
rect 2586 2688 2590 2691
rect 2602 2688 2737 2691
rect 1926 2682 1929 2688
rect 2398 2682 2401 2688
rect 2734 2682 2737 2688
rect 3030 2688 3086 2691
rect 3106 2688 3193 2691
rect 3266 2688 3286 2691
rect 3706 2688 3806 2691
rect 4034 2688 4262 2691
rect 4322 2688 4326 2691
rect 3030 2682 3033 2688
rect 74 2678 222 2681
rect 266 2678 318 2681
rect 322 2678 382 2681
rect 386 2678 438 2681
rect 850 2678 942 2681
rect 1402 2678 1478 2681
rect 1650 2678 1734 2681
rect 1770 2678 1926 2681
rect 2058 2678 2177 2681
rect 2250 2678 2254 2681
rect 2370 2678 2382 2681
rect 2538 2678 2654 2681
rect 2658 2678 2678 2681
rect 3086 2681 3089 2688
rect 3190 2682 3193 2688
rect 3430 2682 3433 2688
rect 3086 2678 3166 2681
rect 3282 2678 3366 2681
rect 3582 2681 3585 2688
rect 3570 2678 3585 2681
rect 3614 2682 3617 2688
rect 3778 2678 3790 2681
rect 3794 2678 3822 2681
rect 3890 2678 3918 2681
rect 3970 2678 3982 2681
rect 3998 2681 4001 2688
rect 3998 2678 4046 2681
rect 4146 2678 4174 2681
rect 4178 2678 4214 2681
rect 146 2668 190 2671
rect 194 2668 238 2671
rect 242 2668 281 2671
rect 298 2668 334 2671
rect 354 2668 598 2671
rect 710 2671 713 2678
rect 710 2668 814 2671
rect 1054 2671 1057 2678
rect 922 2668 1057 2671
rect 1218 2668 1238 2671
rect 1242 2668 1246 2671
rect 1334 2671 1337 2678
rect 1334 2668 1454 2671
rect 1526 2671 1529 2678
rect 1542 2672 1545 2678
rect 2046 2672 2049 2678
rect 1526 2668 1534 2671
rect 1658 2668 1662 2671
rect 1874 2668 1910 2671
rect 2146 2668 2166 2671
rect 2174 2671 2177 2678
rect 2174 2668 2305 2671
rect 2362 2668 2414 2671
rect 2418 2668 2470 2671
rect 2474 2668 2582 2671
rect 2714 2668 2718 2671
rect 2746 2668 2750 2671
rect 2946 2668 2950 2671
rect 3002 2668 3006 2671
rect 3014 2671 3017 2678
rect 3014 2668 3030 2671
rect 3034 2668 3062 2671
rect 3098 2668 3110 2671
rect 3170 2668 3278 2671
rect 3282 2668 3310 2671
rect 3414 2668 3561 2671
rect 3586 2668 3614 2671
rect 3770 2668 3838 2671
rect 4034 2668 4038 2671
rect 4106 2668 4145 2671
rect 4186 2668 4206 2671
rect 4390 2671 4393 2678
rect 4282 2668 4393 2671
rect 278 2662 281 2668
rect 218 2658 254 2661
rect 282 2658 358 2661
rect 378 2658 502 2661
rect 530 2658 534 2661
rect 554 2658 574 2661
rect 674 2658 726 2661
rect 730 2658 1350 2661
rect 1478 2661 1481 2668
rect 2302 2662 2305 2668
rect 2766 2662 2769 2668
rect 3414 2662 3417 2668
rect 3558 2662 3561 2668
rect 1394 2658 1481 2661
rect 1890 2658 1902 2661
rect 2050 2658 2134 2661
rect 2138 2658 2150 2661
rect 2154 2658 2190 2661
rect 2234 2658 2270 2661
rect 2322 2658 2334 2661
rect 2386 2658 2414 2661
rect 2466 2658 2638 2661
rect 2642 2658 2742 2661
rect 2922 2658 3022 2661
rect 3074 2658 3118 2661
rect 3162 2658 3166 2661
rect 3202 2658 3214 2661
rect 3218 2658 3326 2661
rect 3738 2658 3742 2661
rect 3894 2661 3897 2668
rect 3874 2658 3897 2661
rect 3938 2658 3950 2661
rect 4142 2661 4145 2668
rect 4142 2658 4233 2661
rect 4290 2658 4305 2661
rect 4314 2658 4342 2661
rect 2350 2652 2353 2658
rect 2750 2652 2753 2658
rect 178 2648 254 2651
rect 258 2648 302 2651
rect 522 2648 537 2651
rect 562 2648 590 2651
rect 626 2648 646 2651
rect 858 2648 894 2651
rect 1210 2648 1214 2651
rect 1546 2648 1630 2651
rect 1854 2648 2206 2651
rect 2210 2648 2342 2651
rect 2370 2648 2630 2651
rect 2642 2648 2670 2651
rect 2690 2648 2742 2651
rect 2794 2648 2798 2651
rect 2802 2648 3054 2651
rect 3138 2648 3150 2651
rect 3154 2648 3198 2651
rect 3202 2648 3214 2651
rect 3218 2648 3294 2651
rect 3546 2648 3574 2651
rect 3674 2648 3734 2651
rect 3774 2651 3777 2658
rect 4134 2652 4137 2658
rect 4230 2652 4233 2658
rect 3738 2648 3777 2651
rect 3914 2648 3926 2651
rect 3962 2648 4006 2651
rect 4010 2648 4046 2651
rect 4106 2648 4110 2651
rect 4146 2648 4150 2651
rect 4290 2648 4294 2651
rect 4302 2651 4305 2658
rect 4302 2648 4342 2651
rect 534 2642 537 2648
rect 1182 2642 1185 2648
rect 1854 2642 1857 2648
rect 418 2638 526 2641
rect 570 2638 574 2641
rect 1306 2638 1854 2641
rect 2146 2638 2158 2641
rect 2194 2638 2294 2641
rect 2298 2638 2326 2641
rect 2330 2638 2454 2641
rect 2458 2638 2486 2641
rect 2674 2638 2702 2641
rect 2746 2638 3062 2641
rect 3090 2638 3110 2641
rect 3178 2638 3230 2641
rect 3242 2638 3262 2641
rect 3538 2638 3854 2641
rect 4130 2638 4158 2641
rect 4166 2641 4169 2648
rect 4162 2638 4169 2641
rect 214 2632 217 2638
rect 242 2628 614 2631
rect 2058 2628 2198 2631
rect 2202 2628 2254 2631
rect 2278 2628 2334 2631
rect 2338 2628 2374 2631
rect 2426 2628 2574 2631
rect 2578 2628 2814 2631
rect 3058 2628 3126 2631
rect 3130 2628 3142 2631
rect 3186 2628 3246 2631
rect 3250 2628 3374 2631
rect 3554 2628 3793 2631
rect 3842 2628 3846 2631
rect 3906 2628 3934 2631
rect 3954 2628 4022 2631
rect 4122 2628 4158 2631
rect 4194 2628 4222 2631
rect 2278 2622 2281 2628
rect 90 2618 662 2621
rect 666 2618 1246 2621
rect 1266 2618 1326 2621
rect 1442 2618 1470 2621
rect 1810 2618 2174 2621
rect 2178 2618 2182 2621
rect 2186 2618 2270 2621
rect 2374 2621 2377 2628
rect 3790 2622 3793 2628
rect 2374 2618 2585 2621
rect 2722 2618 2750 2621
rect 2818 2618 2822 2621
rect 2842 2618 3182 2621
rect 3522 2618 3606 2621
rect 3634 2618 3766 2621
rect 3770 2618 3774 2621
rect 3794 2618 3998 2621
rect 4090 2618 4350 2621
rect 426 2608 486 2611
rect 546 2608 638 2611
rect 1074 2608 1150 2611
rect 1586 2608 1654 2611
rect 1658 2608 1694 2611
rect 1698 2608 1766 2611
rect 1826 2608 2406 2611
rect 2410 2608 2414 2611
rect 2498 2608 2502 2611
rect 2582 2611 2585 2618
rect 2582 2608 2854 2611
rect 2922 2608 3110 2611
rect 3642 2608 3846 2611
rect 3850 2608 4022 2611
rect 4082 2608 4206 2611
rect 392 2603 394 2607
rect 398 2603 401 2607
rect 406 2603 408 2607
rect 1416 2603 1418 2607
rect 1422 2603 1425 2607
rect 1430 2603 1432 2607
rect 2440 2603 2442 2607
rect 2446 2603 2449 2607
rect 2454 2603 2456 2607
rect 3472 2603 3474 2607
rect 3478 2603 3481 2607
rect 3486 2603 3488 2607
rect 490 2598 550 2601
rect 610 2598 878 2601
rect 1050 2598 1126 2601
rect 1194 2598 1198 2601
rect 1994 2598 2046 2601
rect 2170 2598 2214 2601
rect 2242 2598 2246 2601
rect 2330 2598 2350 2601
rect 2514 2598 2718 2601
rect 2978 2598 3446 2601
rect 3690 2598 3694 2601
rect 3858 2598 3966 2601
rect 3970 2598 4150 2601
rect 38 2592 41 2598
rect 94 2592 97 2598
rect 266 2588 270 2591
rect 1114 2588 1246 2591
rect 1386 2588 1854 2591
rect 1858 2588 2070 2591
rect 2242 2588 2326 2591
rect 2490 2588 2886 2591
rect 4010 2588 4038 2591
rect 4042 2588 4142 2591
rect 506 2578 510 2581
rect 594 2578 598 2581
rect 790 2581 793 2588
rect 790 2578 1390 2581
rect 1394 2578 1542 2581
rect 1786 2578 1894 2581
rect 1898 2578 2398 2581
rect 2402 2578 2726 2581
rect 2730 2578 2790 2581
rect 2826 2578 3054 2581
rect 3090 2578 3310 2581
rect 3346 2578 3558 2581
rect 3610 2578 3662 2581
rect 3666 2578 3854 2581
rect 3886 2581 3889 2588
rect 3886 2578 4014 2581
rect 4042 2578 4246 2581
rect 4250 2578 4270 2581
rect 34 2568 214 2571
rect 514 2568 526 2571
rect 594 2568 630 2571
rect 754 2568 966 2571
rect 970 2568 1614 2571
rect 1754 2568 2214 2571
rect 2346 2568 2486 2571
rect 2546 2568 2558 2571
rect 2634 2568 3150 2571
rect 3330 2568 4006 2571
rect 4014 2571 4017 2578
rect 4014 2568 4078 2571
rect 4138 2568 4214 2571
rect 114 2558 118 2561
rect 202 2558 230 2561
rect 474 2558 649 2561
rect 666 2558 830 2561
rect 1522 2558 1814 2561
rect 1834 2558 1894 2561
rect 1946 2558 2014 2561
rect 2082 2558 2094 2561
rect 2114 2558 2174 2561
rect 2274 2558 2278 2561
rect 2426 2558 2454 2561
rect 2498 2558 2502 2561
rect 2594 2558 2718 2561
rect 2938 2558 3030 2561
rect 3250 2558 3254 2561
rect 3586 2558 3630 2561
rect 3634 2558 3646 2561
rect 3698 2558 3718 2561
rect 3770 2558 3814 2561
rect 3978 2558 4054 2561
rect 4058 2558 4062 2561
rect 4170 2558 4310 2561
rect 4370 2558 4374 2561
rect -26 2551 -22 2552
rect -26 2548 6 2551
rect 210 2548 246 2551
rect 602 2548 606 2551
rect 646 2551 649 2558
rect 646 2548 726 2551
rect 730 2548 758 2551
rect 834 2548 862 2551
rect 1102 2551 1105 2558
rect 1102 2548 1118 2551
rect 1122 2548 1278 2551
rect 1334 2551 1337 2558
rect 1290 2548 1337 2551
rect 1434 2548 1614 2551
rect 1754 2548 1758 2551
rect 1778 2548 1838 2551
rect 1894 2551 1897 2558
rect 1882 2548 1897 2551
rect 1970 2548 2078 2551
rect 2082 2548 2134 2551
rect 2162 2548 2230 2551
rect 2290 2548 2366 2551
rect 2506 2548 2646 2551
rect 2650 2548 2654 2551
rect 2770 2548 2774 2551
rect 2778 2548 2806 2551
rect 2850 2548 2910 2551
rect 3154 2548 3230 2551
rect 3234 2548 3238 2551
rect 3266 2548 3270 2551
rect 3330 2548 3462 2551
rect 3594 2548 3598 2551
rect 3778 2548 3782 2551
rect 3786 2548 3806 2551
rect 3810 2548 3918 2551
rect 3922 2548 4070 2551
rect 4074 2548 4134 2551
rect 4146 2548 4230 2551
rect 118 2541 121 2548
rect 90 2538 121 2541
rect 154 2538 174 2541
rect 194 2538 214 2541
rect 274 2538 478 2541
rect 490 2538 494 2541
rect 514 2538 518 2541
rect 546 2538 590 2541
rect 842 2538 870 2541
rect 950 2541 953 2548
rect 1094 2541 1097 2548
rect 950 2538 1097 2541
rect 1138 2538 1574 2541
rect 1578 2538 1782 2541
rect 1810 2538 1910 2541
rect 1914 2538 1918 2541
rect 2002 2538 2006 2541
rect 2026 2538 2054 2541
rect 2066 2538 2070 2541
rect 2154 2538 2262 2541
rect 2282 2538 2318 2541
rect 2322 2538 2326 2541
rect 2338 2538 2422 2541
rect 2538 2538 2542 2541
rect 2554 2538 2606 2541
rect 2966 2541 2969 2548
rect 2946 2538 2969 2541
rect 3006 2542 3009 2548
rect 3146 2538 3158 2541
rect 3194 2538 3230 2541
rect 3306 2538 3342 2541
rect 3618 2538 3686 2541
rect 3714 2538 3718 2541
rect 3762 2538 3766 2541
rect 3834 2538 3838 2541
rect 3850 2538 3950 2541
rect 4018 2538 4030 2541
rect 4062 2538 4129 2541
rect 4146 2538 4150 2541
rect 4154 2538 4190 2541
rect 4318 2541 4321 2548
rect 4314 2538 4321 2541
rect 26 2528 241 2531
rect 434 2528 486 2531
rect 490 2528 494 2531
rect 570 2528 582 2531
rect 650 2528 662 2531
rect 1242 2528 1294 2531
rect 1506 2528 1510 2531
rect 1602 2528 1630 2531
rect 1634 2528 1673 2531
rect 1770 2528 1854 2531
rect 1870 2528 2038 2531
rect 2042 2528 2070 2531
rect 2098 2528 2102 2531
rect 2178 2528 2198 2531
rect 2226 2528 2262 2531
rect 2266 2528 2270 2531
rect 2298 2528 2302 2531
rect 2314 2528 2342 2531
rect 2426 2528 2430 2531
rect 2554 2528 2598 2531
rect 2602 2528 2622 2531
rect 2658 2528 2662 2531
rect 2794 2528 2910 2531
rect 2950 2528 2974 2531
rect 3166 2531 3169 2538
rect 4062 2532 4065 2538
rect 4126 2532 4129 2538
rect 3166 2528 3206 2531
rect 3258 2528 3278 2531
rect 3298 2528 3334 2531
rect 3394 2528 3550 2531
rect 3610 2528 3654 2531
rect 3674 2528 3758 2531
rect 3762 2528 3774 2531
rect 3842 2528 3870 2531
rect 3874 2528 3894 2531
rect 3946 2528 3966 2531
rect 4002 2528 4022 2531
rect 4298 2528 4318 2531
rect 4362 2528 4390 2531
rect 238 2521 241 2528
rect 238 2518 1078 2521
rect 1142 2521 1145 2528
rect 1670 2522 1673 2528
rect 1870 2522 1873 2528
rect 2350 2522 2353 2528
rect 2950 2522 2953 2528
rect 3838 2522 3841 2528
rect 1142 2518 1238 2521
rect 1554 2518 1558 2521
rect 1562 2518 1665 2521
rect 1954 2518 2030 2521
rect 2034 2518 2158 2521
rect 2170 2518 2222 2521
rect 2258 2518 2334 2521
rect 2370 2518 2462 2521
rect 2546 2518 2574 2521
rect 2602 2518 2670 2521
rect 2674 2518 2686 2521
rect 2698 2518 2702 2521
rect 3062 2518 3102 2521
rect 3106 2518 3214 2521
rect 3226 2518 3286 2521
rect 3322 2518 3358 2521
rect 3506 2518 3566 2521
rect 3618 2518 3622 2521
rect 3858 2518 3950 2521
rect 3954 2518 4086 2521
rect 234 2508 390 2511
rect 394 2508 454 2511
rect 490 2508 542 2511
rect 554 2508 566 2511
rect 578 2508 606 2511
rect 970 2508 1518 2511
rect 1634 2508 1654 2511
rect 1662 2511 1665 2518
rect 3062 2512 3065 2518
rect 1662 2508 1814 2511
rect 2082 2508 2134 2511
rect 2258 2508 2262 2511
rect 2298 2508 2478 2511
rect 2502 2508 2614 2511
rect 2618 2508 2662 2511
rect 2810 2508 2902 2511
rect 2938 2508 2942 2511
rect 3218 2508 3566 2511
rect 3602 2508 3726 2511
rect 3778 2508 3790 2511
rect 3898 2508 3966 2511
rect 896 2503 898 2507
rect 902 2503 905 2507
rect 910 2503 912 2507
rect 1928 2503 1930 2507
rect 1934 2503 1937 2507
rect 1942 2503 1944 2507
rect 74 2498 110 2501
rect 130 2498 166 2501
rect 178 2498 214 2501
rect 338 2498 358 2501
rect 362 2498 790 2501
rect 1042 2498 1150 2501
rect 1154 2498 1438 2501
rect 1450 2498 1790 2501
rect 1802 2498 1918 2501
rect 1962 2498 2006 2501
rect 2010 2498 2014 2501
rect 2018 2498 2126 2501
rect 2130 2498 2142 2501
rect 2178 2498 2310 2501
rect 2502 2501 2505 2508
rect 2952 2503 2954 2507
rect 2958 2503 2961 2507
rect 2966 2503 2968 2507
rect 3976 2503 3978 2507
rect 3982 2503 3985 2507
rect 3990 2503 3992 2507
rect 2386 2498 2505 2501
rect 2514 2498 2598 2501
rect 2602 2498 2710 2501
rect 2714 2498 2774 2501
rect 2778 2498 2945 2501
rect 3130 2498 3246 2501
rect 3282 2498 3318 2501
rect 3418 2498 3662 2501
rect 3666 2498 3742 2501
rect 3746 2498 3846 2501
rect 3850 2498 3969 2501
rect 190 2488 294 2491
rect 298 2488 382 2491
rect 578 2488 582 2491
rect 626 2488 638 2491
rect 642 2488 814 2491
rect 930 2488 1222 2491
rect 1226 2488 1230 2491
rect 1242 2488 1270 2491
rect 1274 2488 1406 2491
rect 1626 2488 1670 2491
rect 1810 2488 1950 2491
rect 2138 2488 2302 2491
rect 2506 2488 2630 2491
rect 2698 2488 2814 2491
rect 2942 2491 2945 2498
rect 3966 2492 3969 2498
rect 2942 2488 2958 2491
rect 3098 2488 3182 2491
rect 3202 2488 3222 2491
rect 3234 2488 3318 2491
rect 3362 2488 3486 2491
rect 3490 2488 3590 2491
rect 3666 2488 3694 2491
rect 3866 2488 3894 2491
rect 3986 2488 4150 2491
rect 4154 2488 4182 2491
rect 4194 2488 4374 2491
rect 86 2482 89 2488
rect 190 2482 193 2488
rect 378 2478 502 2481
rect 594 2478 646 2481
rect 926 2481 929 2488
rect 762 2478 929 2481
rect 970 2478 990 2481
rect 994 2478 1006 2481
rect 1010 2478 1086 2481
rect 1218 2478 1286 2481
rect 1394 2478 1438 2481
rect 1462 2481 1465 2488
rect 1694 2482 1697 2488
rect 1442 2478 1465 2481
rect 1682 2478 1686 2481
rect 1706 2478 1718 2481
rect 1734 2478 1737 2488
rect 1870 2482 1873 2488
rect 1882 2478 1990 2481
rect 2038 2481 2041 2488
rect 2010 2478 2041 2481
rect 2090 2478 2398 2481
rect 2402 2478 2574 2481
rect 2610 2478 2630 2481
rect 2642 2478 2734 2481
rect 3086 2481 3089 2488
rect 2930 2478 3089 2481
rect 3114 2478 3166 2481
rect 3194 2478 3278 2481
rect 3282 2478 3494 2481
rect 3530 2478 3534 2481
rect 3546 2478 3614 2481
rect 3658 2478 3710 2481
rect 3782 2481 3785 2488
rect 3714 2478 3785 2481
rect 3914 2478 3918 2481
rect 3966 2481 3969 2488
rect 3966 2478 4022 2481
rect 4082 2478 4134 2481
rect 4234 2478 4238 2481
rect 310 2471 313 2478
rect 242 2468 313 2471
rect 550 2471 553 2478
rect 1046 2472 1049 2478
rect 550 2468 630 2471
rect 658 2468 1014 2471
rect 1058 2468 1137 2471
rect 1282 2468 1366 2471
rect 1370 2468 1425 2471
rect 1434 2468 1481 2471
rect 1522 2468 1598 2471
rect 1634 2468 1646 2471
rect 1674 2468 1710 2471
rect 1754 2468 1854 2471
rect 1874 2468 1886 2471
rect 1938 2468 2054 2471
rect 2058 2468 2094 2471
rect 2250 2468 2262 2471
rect 2490 2468 2518 2471
rect 2522 2468 2558 2471
rect 2586 2468 2606 2471
rect 2646 2468 2678 2471
rect 2698 2468 2702 2471
rect 2746 2468 2750 2471
rect 2754 2468 2798 2471
rect 2818 2468 2982 2471
rect 3002 2468 3006 2471
rect 3082 2468 3134 2471
rect 3162 2468 3190 2471
rect 3202 2468 3206 2471
rect 3242 2468 3254 2471
rect 3298 2468 3318 2471
rect 3322 2468 3326 2471
rect 3362 2468 3366 2471
rect 3386 2468 3430 2471
rect 3450 2468 3494 2471
rect 3538 2468 3542 2471
rect 3546 2468 3622 2471
rect 3626 2468 3686 2471
rect 3698 2468 3718 2471
rect 3866 2468 4078 2471
rect 4178 2468 4222 2471
rect 4306 2468 4326 2471
rect 4330 2468 4358 2471
rect 1134 2462 1137 2468
rect 298 2458 414 2461
rect 546 2458 614 2461
rect 746 2458 750 2461
rect 1330 2458 1358 2461
rect 1370 2458 1374 2461
rect 1422 2461 1425 2468
rect 1422 2458 1470 2461
rect 1478 2461 1481 2468
rect 2646 2462 2649 2468
rect 1478 2458 1654 2461
rect 1658 2458 1662 2461
rect 1690 2458 1830 2461
rect 1834 2458 1838 2461
rect 1866 2458 1894 2461
rect 1962 2458 1974 2461
rect 2010 2458 2025 2461
rect 2050 2458 2054 2461
rect 2074 2458 2118 2461
rect 2122 2458 2326 2461
rect 2330 2458 2358 2461
rect 2370 2458 2374 2461
rect 2490 2458 2590 2461
rect 2738 2458 2750 2461
rect 2818 2458 2870 2461
rect 2914 2458 3038 2461
rect 3042 2458 3246 2461
rect 3274 2458 3302 2461
rect 3306 2458 3310 2461
rect 3322 2458 3342 2461
rect 3362 2458 3422 2461
rect 3522 2458 3526 2461
rect 3538 2458 3630 2461
rect 3666 2458 3670 2461
rect 3778 2458 3814 2461
rect 3938 2458 3982 2461
rect 4090 2458 4110 2461
rect 4138 2458 4174 2461
rect 4178 2458 4270 2461
rect 4298 2458 4350 2461
rect 1070 2452 1073 2458
rect 2022 2452 2025 2458
rect 2782 2452 2785 2458
rect 34 2450 38 2451
rect 30 2448 38 2450
rect 42 2448 366 2451
rect 370 2448 422 2451
rect 506 2448 510 2451
rect 618 2448 622 2451
rect 1098 2448 1342 2451
rect 1346 2448 1350 2451
rect 1378 2448 1486 2451
rect 1506 2448 1542 2451
rect 1546 2448 1582 2451
rect 1618 2448 1750 2451
rect 1754 2448 1806 2451
rect 1978 2448 1982 2451
rect 2082 2448 2086 2451
rect 2218 2448 2262 2451
rect 2338 2448 2390 2451
rect 2410 2448 2446 2451
rect 2490 2448 2614 2451
rect 2754 2448 2758 2451
rect 2858 2448 2918 2451
rect 3066 2448 3070 2451
rect 3146 2448 3166 2451
rect 3194 2448 3278 2451
rect 3334 2448 3342 2451
rect 3346 2448 3462 2451
rect 3546 2448 3566 2451
rect 4070 2451 4073 2458
rect 4026 2448 4073 2451
rect 4218 2448 4294 2451
rect 4338 2448 4382 2451
rect 3134 2442 3137 2448
rect 418 2438 726 2441
rect 1066 2438 1270 2441
rect 1306 2438 1366 2441
rect 1370 2438 1518 2441
rect 1522 2438 1566 2441
rect 1586 2438 1630 2441
rect 1650 2438 1654 2441
rect 1746 2438 1774 2441
rect 1906 2438 2038 2441
rect 2042 2438 2070 2441
rect 2354 2438 2358 2441
rect 2418 2438 2502 2441
rect 2506 2438 2798 2441
rect 2826 2438 2894 2441
rect 2898 2438 3118 2441
rect 3178 2438 3262 2441
rect 3274 2438 3846 2441
rect 3850 2438 3926 2441
rect 3930 2438 3998 2441
rect 4002 2438 4094 2441
rect 4158 2441 4161 2448
rect 4158 2438 4318 2441
rect 4322 2438 4342 2441
rect 1550 2432 1553 2438
rect 1798 2432 1801 2438
rect 482 2428 590 2431
rect 1322 2428 1494 2431
rect 1642 2428 1662 2431
rect 1714 2428 1742 2431
rect 1826 2428 2110 2431
rect 2170 2428 2494 2431
rect 2498 2428 2686 2431
rect 2754 2428 2758 2431
rect 2770 2428 3150 2431
rect 3170 2428 3494 2431
rect 3658 2428 3662 2431
rect 3730 2428 3798 2431
rect 3802 2428 3998 2431
rect 442 2418 526 2421
rect 530 2418 574 2421
rect 578 2418 622 2421
rect 730 2418 1206 2421
rect 1338 2418 1382 2421
rect 1502 2421 1505 2428
rect 3606 2422 3609 2428
rect 1458 2418 1505 2421
rect 1586 2418 1830 2421
rect 1842 2418 2030 2421
rect 2034 2418 2230 2421
rect 2298 2418 2310 2421
rect 2322 2418 2566 2421
rect 2570 2418 2846 2421
rect 2850 2418 2950 2421
rect 2954 2418 2998 2421
rect 3002 2418 3142 2421
rect 3178 2418 3398 2421
rect 3402 2418 3406 2421
rect 4162 2418 4174 2421
rect 498 2408 558 2411
rect 562 2408 1150 2411
rect 1154 2408 1230 2411
rect 1442 2408 1510 2411
rect 1530 2408 1638 2411
rect 1642 2408 1686 2411
rect 1754 2408 1998 2411
rect 2002 2408 2006 2411
rect 2018 2408 2350 2411
rect 2354 2408 2430 2411
rect 2650 2408 2790 2411
rect 2794 2408 2878 2411
rect 3034 2408 3310 2411
rect 3794 2408 4262 2411
rect 4266 2408 4286 2411
rect 392 2403 394 2407
rect 398 2403 401 2407
rect 406 2403 408 2407
rect 1416 2403 1418 2407
rect 1422 2403 1425 2407
rect 1430 2403 1432 2407
rect 890 2398 910 2401
rect 1186 2398 1214 2401
rect 1354 2398 1398 2401
rect 1526 2401 1529 2408
rect 2440 2403 2442 2407
rect 2446 2403 2449 2407
rect 2454 2403 2456 2407
rect 3472 2403 3474 2407
rect 3478 2403 3481 2407
rect 3486 2403 3488 2407
rect 1466 2398 1529 2401
rect 1682 2398 1758 2401
rect 1850 2398 1910 2401
rect 1914 2398 2422 2401
rect 2426 2398 2430 2401
rect 2754 2398 2838 2401
rect 2978 2398 3465 2401
rect 4242 2398 4254 2401
rect 1402 2388 1406 2391
rect 1410 2388 1478 2391
rect 1530 2388 1702 2391
rect 1830 2391 1833 2398
rect 1738 2388 1833 2391
rect 1954 2388 1982 2391
rect 1986 2388 2126 2391
rect 2130 2388 2158 2391
rect 2282 2388 2678 2391
rect 2778 2388 2822 2391
rect 2842 2388 3406 2391
rect 3462 2391 3465 2398
rect 3462 2388 3734 2391
rect 4202 2388 4214 2391
rect 1810 2378 1814 2381
rect 1818 2378 2062 2381
rect 2082 2378 2246 2381
rect 2250 2378 2406 2381
rect 2418 2378 2654 2381
rect 2874 2378 3014 2381
rect 3026 2378 3038 2381
rect 3050 2378 3166 2381
rect 3618 2378 3630 2381
rect 3826 2378 4062 2381
rect 866 2368 1078 2371
rect 1126 2371 1129 2378
rect 1098 2368 1129 2371
rect 1134 2372 1137 2378
rect 1146 2368 1158 2371
rect 1186 2368 1310 2371
rect 1454 2368 1750 2371
rect 1778 2368 1806 2371
rect 1914 2368 1958 2371
rect 1978 2368 1990 2371
rect 2058 2368 2118 2371
rect 2146 2368 2206 2371
rect 2226 2368 2302 2371
rect 2546 2368 2566 2371
rect 2578 2368 2582 2371
rect 2610 2368 2630 2371
rect 2634 2368 2641 2371
rect 2650 2368 2654 2371
rect 2666 2368 2766 2371
rect 2806 2371 2809 2378
rect 2806 2368 2910 2371
rect 2914 2368 3014 2371
rect 3018 2368 3094 2371
rect 3182 2371 3185 2378
rect 3182 2368 3238 2371
rect 3258 2368 3550 2371
rect 3586 2368 3798 2371
rect 3906 2368 3926 2371
rect 3970 2368 4054 2371
rect 4106 2368 4118 2371
rect 1454 2362 1457 2368
rect 362 2358 670 2361
rect 1082 2358 1105 2361
rect 1122 2358 1342 2361
rect 1658 2358 1686 2361
rect 1714 2358 1750 2361
rect 1834 2358 1950 2361
rect 1978 2358 2150 2361
rect 2178 2358 2241 2361
rect 2482 2358 2486 2361
rect 2522 2358 2774 2361
rect 2794 2358 2798 2361
rect 2802 2358 2862 2361
rect 2882 2358 2902 2361
rect 2930 2358 2974 2361
rect 3010 2358 3134 2361
rect 3162 2358 3166 2361
rect 3170 2358 3190 2361
rect 3298 2358 3326 2361
rect 3338 2358 3470 2361
rect 3574 2358 3582 2361
rect 3586 2358 3598 2361
rect 3826 2358 3846 2361
rect 3850 2358 3894 2361
rect 4026 2358 4134 2361
rect 4150 2361 4153 2368
rect 4182 2361 4185 2368
rect 4358 2362 4361 2368
rect 4374 2362 4377 2368
rect 4150 2358 4185 2361
rect 4226 2358 4230 2361
rect 1102 2352 1105 2358
rect 1790 2352 1793 2358
rect 194 2348 222 2351
rect 226 2348 286 2351
rect 618 2348 726 2351
rect 842 2348 878 2351
rect 1106 2348 1158 2351
rect 1162 2348 1318 2351
rect 1322 2348 1342 2351
rect 1386 2348 1390 2351
rect 1498 2348 1534 2351
rect 1666 2348 1686 2351
rect 1690 2348 1718 2351
rect 1762 2348 1774 2351
rect 1814 2351 1817 2358
rect 2238 2352 2241 2358
rect 3902 2352 3905 2358
rect 1802 2348 1817 2351
rect 1858 2348 1942 2351
rect 1946 2348 2038 2351
rect 2082 2348 2118 2351
rect 2122 2348 2166 2351
rect 2186 2348 2190 2351
rect 2210 2348 2222 2351
rect 2330 2348 2342 2351
rect 2362 2348 2462 2351
rect 2482 2348 2590 2351
rect 2746 2348 2774 2351
rect 2778 2348 2814 2351
rect 2850 2348 2878 2351
rect 2882 2348 2998 2351
rect 3066 2348 3081 2351
rect 134 2341 137 2348
rect 2038 2342 2041 2348
rect 3078 2342 3081 2348
rect 3114 2348 3174 2351
rect 3202 2348 3222 2351
rect 3274 2348 3302 2351
rect 3314 2348 3358 2351
rect 3362 2348 3406 2351
rect 3522 2348 3630 2351
rect 4010 2348 4014 2351
rect 4122 2348 4198 2351
rect 4202 2348 4254 2351
rect 4342 2351 4345 2358
rect 4382 2352 4385 2358
rect 4274 2348 4366 2351
rect 3086 2342 3089 2348
rect 34 2338 137 2341
rect 178 2338 214 2341
rect 218 2338 430 2341
rect 434 2338 470 2341
rect 934 2338 1006 2341
rect 1058 2338 1062 2341
rect 1066 2338 1142 2341
rect 1210 2338 1270 2341
rect 1322 2338 1358 2341
rect 1386 2338 1390 2341
rect 1402 2338 1406 2341
rect 1522 2338 1542 2341
rect 1546 2338 1630 2341
rect 1658 2338 1670 2341
rect 1674 2338 1694 2341
rect 1722 2338 1830 2341
rect 1858 2338 1862 2341
rect 1890 2338 1894 2341
rect 1902 2338 1966 2341
rect 1994 2338 1998 2341
rect 2074 2338 2094 2341
rect 2106 2338 2126 2341
rect 2218 2338 2278 2341
rect 2394 2338 2454 2341
rect 2466 2338 2494 2341
rect 2498 2338 2518 2341
rect 2530 2338 2574 2341
rect 2634 2338 2638 2341
rect 2674 2338 2678 2341
rect 2682 2338 2750 2341
rect 2794 2338 2833 2341
rect 2842 2338 2886 2341
rect 2898 2338 2934 2341
rect 2994 2338 3022 2341
rect 3138 2338 3230 2341
rect 3258 2338 3278 2341
rect 3306 2338 3342 2341
rect 3554 2338 3558 2341
rect 3570 2338 3574 2341
rect 3818 2338 3822 2341
rect 3866 2338 3870 2341
rect 4202 2338 4206 2341
rect 4314 2338 4318 2341
rect 4322 2338 4326 2341
rect 90 2328 121 2331
rect 346 2328 377 2331
rect 566 2331 569 2338
rect 386 2328 569 2331
rect 578 2328 662 2331
rect 766 2331 769 2338
rect 666 2328 769 2331
rect 934 2332 937 2338
rect 962 2328 1014 2331
rect 1018 2328 1030 2331
rect 1098 2328 1142 2331
rect 1502 2331 1505 2338
rect 1482 2328 1505 2331
rect 1610 2328 1614 2331
rect 1650 2328 1758 2331
rect 1770 2328 1814 2331
rect 1818 2328 1822 2331
rect 1902 2331 1905 2338
rect 2342 2332 2345 2338
rect 1874 2328 1905 2331
rect 1970 2328 2062 2331
rect 2090 2328 2094 2331
rect 2138 2328 2230 2331
rect 2258 2328 2342 2331
rect 2402 2328 2534 2331
rect 2558 2328 2566 2331
rect 2570 2328 2678 2331
rect 2690 2328 2694 2331
rect 2702 2328 2710 2331
rect 2714 2328 2766 2331
rect 2770 2328 2822 2331
rect 2830 2331 2833 2338
rect 3358 2332 3361 2338
rect 2830 2328 2854 2331
rect 2978 2328 3006 2331
rect 3034 2328 3070 2331
rect 3162 2328 3182 2331
rect 3202 2328 3206 2331
rect 3234 2328 3270 2331
rect 3282 2328 3334 2331
rect 3626 2328 3686 2331
rect 3858 2328 3862 2331
rect 3898 2328 4006 2331
rect 4034 2328 4222 2331
rect 118 2322 121 2328
rect 122 2318 366 2321
rect 374 2321 377 2328
rect 1254 2322 1257 2328
rect 374 2318 662 2321
rect 698 2318 710 2321
rect 714 2318 726 2321
rect 1090 2318 1158 2321
rect 1162 2318 1174 2321
rect 1606 2321 1609 2328
rect 1458 2318 1609 2321
rect 1622 2322 1625 2328
rect 1666 2318 2086 2321
rect 2090 2318 2254 2321
rect 2346 2318 2446 2321
rect 2578 2318 2814 2321
rect 2818 2318 2822 2321
rect 2834 2318 3078 2321
rect 3082 2318 3206 2321
rect 3214 2321 3217 2328
rect 3214 2318 3230 2321
rect 3338 2318 3366 2321
rect 3506 2318 3590 2321
rect 3594 2318 3614 2321
rect 3898 2318 3934 2321
rect 3954 2318 4038 2321
rect 4074 2318 4222 2321
rect 4354 2318 4358 2321
rect -26 2311 -22 2312
rect -26 2308 22 2311
rect 554 2308 694 2311
rect 746 2308 750 2311
rect 986 2308 1046 2311
rect 1082 2308 1110 2311
rect 1114 2308 1318 2311
rect 1498 2308 1670 2311
rect 1698 2308 1758 2311
rect 1778 2308 1846 2311
rect 1866 2308 1870 2311
rect 1970 2308 2022 2311
rect 2042 2308 2134 2311
rect 2146 2308 2470 2311
rect 2474 2308 2550 2311
rect 2562 2308 2750 2311
rect 3194 2308 3262 2311
rect 3274 2308 3302 2311
rect 3346 2308 3766 2311
rect 4218 2308 4254 2311
rect 4258 2308 4286 2311
rect 4354 2308 4374 2311
rect 896 2303 898 2307
rect 902 2303 905 2307
rect 910 2303 912 2307
rect 1928 2303 1930 2307
rect 1934 2303 1937 2307
rect 1942 2303 1944 2307
rect 2952 2303 2954 2307
rect 2958 2303 2961 2307
rect 2966 2303 2968 2307
rect 3976 2303 3978 2307
rect 3982 2303 3985 2307
rect 3990 2303 3992 2307
rect 538 2298 566 2301
rect 746 2298 790 2301
rect 794 2298 822 2301
rect 938 2298 1094 2301
rect 1218 2298 1246 2301
rect 1250 2298 1390 2301
rect 1442 2298 1446 2301
rect 1682 2298 1710 2301
rect 1754 2298 1862 2301
rect 1882 2298 1910 2301
rect 1986 2298 1990 2301
rect 2034 2298 2094 2301
rect 2098 2298 2182 2301
rect 2266 2298 2366 2301
rect 2370 2298 2614 2301
rect 3210 2298 3358 2301
rect 3362 2298 3398 2301
rect 3410 2298 3590 2301
rect 3706 2298 3886 2301
rect 3922 2298 3942 2301
rect 4066 2298 4310 2301
rect 4314 2298 4350 2301
rect -26 2291 -22 2292
rect -26 2288 65 2291
rect 62 2282 65 2288
rect 194 2288 1046 2291
rect 1058 2288 1510 2291
rect 1602 2288 1662 2291
rect 1682 2288 3422 2291
rect 3434 2288 3454 2291
rect 3458 2288 3513 2291
rect 3610 2288 3678 2291
rect 4090 2288 4094 2291
rect 4154 2288 4166 2291
rect 4266 2288 4318 2291
rect 174 2281 177 2288
rect 170 2278 262 2281
rect 674 2278 822 2281
rect 826 2278 886 2281
rect 906 2278 950 2281
rect 954 2278 958 2281
rect 978 2278 1022 2281
rect 1026 2278 1030 2281
rect 1322 2278 1334 2281
rect 1442 2278 1449 2281
rect 1594 2278 1606 2281
rect 1610 2278 1617 2281
rect 1642 2278 1646 2281
rect 1666 2278 1670 2281
rect 1698 2278 1702 2281
rect 1722 2278 1726 2281
rect 1778 2278 1806 2281
rect 1842 2278 1862 2281
rect 1866 2278 1902 2281
rect 1906 2278 1974 2281
rect 1978 2278 2078 2281
rect 2082 2278 2102 2281
rect 2274 2278 2398 2281
rect 2458 2278 2494 2281
rect 2506 2278 2662 2281
rect 2734 2278 2766 2281
rect 3186 2278 3414 2281
rect 3434 2278 3502 2281
rect 3510 2281 3513 2288
rect 3510 2278 3694 2281
rect 3858 2278 3862 2281
rect 3914 2278 3918 2281
rect 3986 2278 3990 2281
rect 4002 2278 4006 2281
rect 4018 2278 4086 2281
rect 4090 2278 4166 2281
rect 4210 2278 4214 2281
rect 4254 2281 4257 2288
rect 4254 2278 4262 2281
rect 4306 2278 4326 2281
rect 4330 2278 4366 2281
rect -26 2271 -22 2272
rect -26 2268 17 2271
rect 34 2268 38 2271
rect 578 2268 606 2271
rect 658 2268 686 2271
rect 690 2268 734 2271
rect 738 2268 766 2271
rect 770 2268 918 2271
rect 922 2268 982 2271
rect 1190 2268 1198 2271
rect 1210 2268 1302 2271
rect 1306 2268 1310 2271
rect 1446 2271 1449 2278
rect 2734 2272 2737 2278
rect 1402 2268 1734 2271
rect 1738 2268 2014 2271
rect 2018 2268 2222 2271
rect 2338 2268 2342 2271
rect 2354 2268 2390 2271
rect 2394 2268 2398 2271
rect 2426 2268 2446 2271
rect 2562 2268 2582 2271
rect 2586 2268 2606 2271
rect 2942 2271 2945 2278
rect 3134 2271 3137 2278
rect 2942 2268 3089 2271
rect 3134 2268 3142 2271
rect 3202 2268 3326 2271
rect 3330 2268 3422 2271
rect 3466 2268 3542 2271
rect 3546 2268 3550 2271
rect 3554 2268 3662 2271
rect 3690 2268 3702 2271
rect 3738 2268 3742 2271
rect 3746 2268 3782 2271
rect 3858 2268 4150 2271
rect 4174 2271 4177 2278
rect 4174 2268 4190 2271
rect 4194 2268 4198 2271
rect 4210 2268 4246 2271
rect 4258 2268 4294 2271
rect 4298 2268 4334 2271
rect 14 2261 17 2268
rect 1190 2262 1193 2268
rect 14 2258 22 2261
rect 426 2258 462 2261
rect 522 2258 654 2261
rect 722 2258 758 2261
rect 762 2258 798 2261
rect 810 2258 814 2261
rect 826 2258 830 2261
rect 842 2258 846 2261
rect 882 2258 926 2261
rect 1034 2258 1038 2261
rect 1122 2258 1126 2261
rect 1522 2258 1606 2261
rect 1674 2258 1734 2261
rect 1762 2258 1854 2261
rect 1858 2258 1870 2261
rect 1906 2258 1998 2261
rect 2002 2258 2006 2261
rect 2018 2258 2030 2261
rect 2138 2258 2142 2261
rect 2322 2258 2342 2261
rect 2378 2258 2574 2261
rect 2594 2258 2758 2261
rect 2810 2258 2854 2261
rect 2858 2258 2886 2261
rect 3002 2258 3006 2261
rect 3010 2258 3078 2261
rect 3086 2261 3089 2268
rect 3086 2258 3230 2261
rect 3258 2258 3334 2261
rect 3370 2258 3374 2261
rect 3394 2258 3398 2261
rect 3410 2258 3454 2261
rect 3458 2258 3550 2261
rect 3554 2258 3561 2261
rect 3570 2258 3582 2261
rect 3594 2258 3646 2261
rect 3710 2261 3713 2268
rect 3650 2258 3750 2261
rect 3754 2258 3782 2261
rect 3826 2258 3838 2261
rect 3946 2258 3998 2261
rect 4026 2258 4038 2261
rect 4058 2258 4238 2261
rect 4242 2258 4262 2261
rect 4290 2258 4294 2261
rect -26 2251 -22 2252
rect 6 2251 9 2258
rect 3294 2252 3297 2258
rect 3350 2252 3353 2258
rect -26 2248 38 2251
rect 714 2248 793 2251
rect 826 2248 878 2251
rect 886 2248 1094 2251
rect 1314 2248 1550 2251
rect 1634 2248 1638 2251
rect 1690 2248 1694 2251
rect 1786 2248 1806 2251
rect 1870 2248 1918 2251
rect 1930 2248 1942 2251
rect 1986 2248 1990 2251
rect 2034 2248 2038 2251
rect 2082 2248 2198 2251
rect 2234 2248 2510 2251
rect 2642 2248 2926 2251
rect 3130 2248 3254 2251
rect 3306 2248 3321 2251
rect 3386 2248 3478 2251
rect 3490 2248 3526 2251
rect 3562 2248 3574 2251
rect 3634 2248 3654 2251
rect 3658 2248 3729 2251
rect 790 2242 793 2248
rect 370 2238 601 2241
rect 850 2238 854 2241
rect 886 2241 889 2248
rect 1782 2242 1785 2248
rect 1870 2242 1873 2248
rect 2014 2242 2017 2248
rect 3318 2242 3321 2248
rect 3726 2242 3729 2248
rect 3938 2248 3950 2251
rect 4130 2248 4142 2251
rect 4146 2248 4182 2251
rect 858 2238 889 2241
rect 954 2238 1326 2241
rect 1570 2238 1686 2241
rect 1818 2238 1865 2241
rect 1886 2238 1902 2241
rect 1906 2238 1918 2241
rect 1954 2238 2006 2241
rect 2386 2238 2486 2241
rect 2546 2238 3030 2241
rect 3034 2238 3246 2241
rect 3330 2238 3529 2241
rect 3610 2238 3718 2241
rect 3838 2241 3841 2248
rect 4062 2242 4065 2248
rect 3818 2238 3841 2241
rect 3882 2238 3886 2241
rect 3890 2238 4030 2241
rect 54 2228 590 2231
rect 598 2231 601 2238
rect 598 2228 774 2231
rect 802 2228 862 2231
rect 1010 2228 1022 2231
rect 1074 2228 1310 2231
rect 1322 2228 1574 2231
rect 1610 2228 1758 2231
rect 1762 2228 1774 2231
rect 1786 2228 1790 2231
rect 1818 2228 1830 2231
rect 1862 2231 1865 2238
rect 1886 2231 1889 2238
rect 3526 2232 3529 2238
rect 1862 2228 1889 2231
rect 1914 2228 1974 2231
rect 1994 2228 2046 2231
rect 2098 2228 2510 2231
rect 2514 2228 2566 2231
rect 2578 2228 2750 2231
rect 2770 2228 3118 2231
rect 3122 2228 3198 2231
rect 3242 2228 3454 2231
rect 3570 2228 3662 2231
rect 3778 2228 3822 2231
rect 3878 2231 3881 2238
rect 3826 2228 3881 2231
rect 3938 2228 4390 2231
rect 54 2222 57 2228
rect 514 2218 518 2221
rect 674 2218 870 2221
rect 966 2221 969 2228
rect 966 2218 974 2221
rect 1018 2218 1038 2221
rect 1282 2218 1286 2221
rect 1450 2218 1518 2221
rect 1546 2218 2030 2221
rect 2034 2218 2406 2221
rect 2546 2218 2638 2221
rect 2642 2218 2646 2221
rect 2826 2218 2838 2221
rect 2842 2218 2846 2221
rect 3306 2218 3702 2221
rect 3910 2218 3918 2221
rect 3922 2218 4014 2221
rect 642 2208 942 2211
rect 946 2208 1046 2211
rect 1178 2208 1182 2211
rect 1362 2208 1382 2211
rect 1538 2208 1606 2211
rect 1610 2208 1678 2211
rect 1698 2208 1886 2211
rect 1890 2208 2286 2211
rect 2626 2208 3230 2211
rect 3242 2208 3334 2211
rect 3498 2208 3558 2211
rect 3562 2208 3758 2211
rect 3762 2208 3846 2211
rect 3850 2208 3910 2211
rect 392 2203 394 2207
rect 398 2203 401 2207
rect 406 2203 408 2207
rect 1416 2203 1418 2207
rect 1422 2203 1425 2207
rect 1430 2203 1432 2207
rect 2440 2203 2442 2207
rect 2446 2203 2449 2207
rect 2454 2203 2456 2207
rect 3472 2203 3474 2207
rect 3478 2203 3481 2207
rect 3486 2203 3488 2207
rect 426 2198 550 2201
rect 554 2198 942 2201
rect 946 2198 1286 2201
rect 1498 2198 1510 2201
rect 1658 2198 2006 2201
rect 2026 2198 2062 2201
rect 2186 2198 2302 2201
rect 2306 2198 2390 2201
rect 2506 2198 2694 2201
rect 2698 2198 2982 2201
rect 3082 2198 3430 2201
rect 3498 2198 3606 2201
rect 3866 2198 3902 2201
rect 3906 2198 3958 2201
rect -26 2191 -22 2192
rect -26 2188 57 2191
rect 258 2188 270 2191
rect 274 2188 318 2191
rect 618 2188 710 2191
rect 718 2188 1158 2191
rect 1162 2188 1390 2191
rect 1394 2188 1630 2191
rect 1666 2188 2214 2191
rect 2322 2188 2358 2191
rect 2370 2188 2718 2191
rect 2882 2188 2910 2191
rect 2962 2188 3174 2191
rect 3274 2188 3425 2191
rect 3522 2188 3593 2191
rect 3850 2188 4022 2191
rect 54 2182 57 2188
rect 618 2178 702 2181
rect 718 2181 721 2188
rect 710 2178 721 2181
rect 746 2178 814 2181
rect 826 2178 846 2181
rect 1186 2178 1398 2181
rect 2278 2181 2281 2188
rect 1626 2178 2081 2181
rect 2278 2178 2318 2181
rect 2322 2178 2326 2181
rect 2370 2178 2478 2181
rect 2482 2178 2526 2181
rect 2530 2178 2550 2181
rect 2730 2178 2894 2181
rect 3230 2181 3233 2188
rect 3422 2182 3425 2188
rect 3590 2182 3593 2188
rect 3230 2178 3262 2181
rect 3282 2178 3286 2181
rect 3378 2178 3414 2181
rect 3778 2178 4134 2181
rect 4150 2181 4153 2188
rect 4150 2178 4214 2181
rect -26 2171 -22 2172
rect 6 2171 9 2178
rect -26 2168 9 2171
rect 710 2171 713 2178
rect 966 2172 969 2178
rect 2078 2172 2081 2178
rect 314 2168 713 2171
rect 718 2168 726 2171
rect 730 2168 734 2171
rect 738 2168 758 2171
rect 762 2168 798 2171
rect 802 2168 830 2171
rect 842 2168 846 2171
rect 874 2168 958 2171
rect 1010 2168 1014 2171
rect 1058 2168 1070 2171
rect 1746 2168 2062 2171
rect 2066 2168 2070 2171
rect 2082 2168 2118 2171
rect 2170 2168 2214 2171
rect 2322 2168 2558 2171
rect 2994 2168 2998 2171
rect 3002 2168 3182 2171
rect 3242 2168 3470 2171
rect 3474 2168 3526 2171
rect 3546 2168 3590 2171
rect 3594 2168 3734 2171
rect 3858 2168 3966 2171
rect 3970 2168 4062 2171
rect -26 2158 30 2161
rect 74 2158 262 2161
rect 642 2158 702 2161
rect 706 2158 998 2161
rect 1002 2158 1110 2161
rect 1114 2158 1150 2161
rect 1382 2161 1385 2168
rect 1322 2158 1385 2161
rect 1434 2158 1438 2161
rect 1686 2161 1689 2168
rect 1686 2158 1729 2161
rect 1738 2158 1758 2161
rect 1770 2158 1806 2161
rect 1834 2158 1966 2161
rect 1978 2158 2030 2161
rect 2034 2158 2038 2161
rect 2058 2158 2150 2161
rect 2218 2158 2366 2161
rect 2410 2158 2414 2161
rect 2578 2158 3158 2161
rect 3162 2158 3286 2161
rect 3290 2158 3510 2161
rect 3682 2158 3702 2161
rect 3738 2158 3758 2161
rect 3762 2158 3774 2161
rect 3802 2158 3806 2161
rect 3954 2158 4062 2161
rect 4074 2158 4078 2161
rect 4166 2161 4169 2168
rect 4166 2158 4190 2161
rect 4230 2161 4233 2168
rect 4230 2158 4262 2161
rect -26 2152 -23 2158
rect -26 2148 -22 2152
rect 26 2148 30 2151
rect 46 2148 54 2151
rect 58 2148 78 2151
rect 202 2148 302 2151
rect 346 2148 766 2151
rect 770 2148 814 2151
rect 842 2148 846 2151
rect 866 2148 926 2151
rect 930 2148 958 2151
rect 962 2148 1382 2151
rect 1518 2148 1614 2151
rect 1618 2148 1670 2151
rect 1674 2148 1705 2151
rect 182 2142 185 2148
rect 630 2138 678 2141
rect 714 2138 758 2141
rect 794 2138 806 2141
rect 818 2138 838 2141
rect 874 2138 878 2141
rect 906 2138 910 2141
rect 922 2138 929 2141
rect 938 2138 942 2141
rect 1018 2138 1078 2141
rect 1098 2138 1118 2141
rect 1306 2138 1310 2141
rect 1518 2141 1521 2148
rect 1702 2142 1705 2148
rect 1726 2151 1729 2158
rect 2198 2152 2201 2158
rect 1726 2148 1798 2151
rect 1906 2148 1910 2151
rect 2010 2148 2046 2151
rect 2050 2148 2062 2151
rect 2298 2148 2302 2151
rect 2450 2148 2486 2151
rect 2490 2148 2497 2151
rect 2570 2148 2654 2151
rect 2674 2148 2678 2151
rect 2682 2148 2734 2151
rect 2842 2148 3166 2151
rect 3202 2148 3206 2151
rect 3218 2148 3246 2151
rect 3250 2148 3257 2151
rect 3290 2148 3294 2151
rect 3354 2148 3358 2151
rect 3362 2148 3414 2151
rect 3418 2148 3542 2151
rect 3566 2151 3569 2158
rect 3566 2148 3638 2151
rect 3642 2148 3718 2151
rect 3778 2148 3782 2151
rect 3906 2148 3998 2151
rect 4046 2148 4054 2151
rect 4098 2148 4102 2151
rect 4162 2148 4174 2151
rect 4202 2148 4238 2151
rect 4354 2148 4366 2151
rect 1370 2138 1521 2141
rect 1650 2138 1678 2141
rect 1718 2141 1721 2148
rect 2822 2142 2825 2148
rect 1718 2138 1774 2141
rect 1850 2138 1934 2141
rect 1954 2138 1990 2141
rect 2002 2138 2006 2141
rect 2050 2138 2110 2141
rect 2118 2138 2126 2141
rect 2130 2138 2177 2141
rect 2258 2138 2262 2141
rect 2266 2138 2286 2141
rect 2330 2138 2334 2141
rect 2354 2138 2534 2141
rect 2578 2138 2582 2141
rect 2658 2138 2686 2141
rect 2902 2138 2910 2141
rect 2914 2138 2942 2141
rect 2946 2138 3238 2141
rect 3258 2138 3318 2141
rect 3346 2138 3374 2141
rect 3426 2138 3462 2141
rect 3546 2138 3697 2141
rect 3706 2138 3710 2141
rect 3730 2138 3734 2141
rect 3754 2138 3806 2141
rect 3814 2138 3838 2141
rect 3970 2138 4102 2141
rect 4130 2138 4150 2141
rect 4154 2138 4222 2141
rect 4278 2141 4281 2148
rect 4278 2138 4382 2141
rect 166 2131 169 2138
rect 166 2128 174 2131
rect 614 2131 617 2138
rect 338 2128 617 2131
rect 630 2132 633 2138
rect 1230 2132 1233 2138
rect 1526 2132 1529 2138
rect 2174 2132 2177 2138
rect 2590 2132 2593 2138
rect 754 2128 766 2131
rect 882 2128 918 2131
rect 1034 2128 1054 2131
rect 1074 2128 1166 2131
rect 1250 2128 1334 2131
rect 1362 2128 1414 2131
rect 1602 2128 1617 2131
rect 1690 2128 1726 2131
rect 1762 2128 1998 2131
rect 2018 2128 2054 2131
rect 2066 2128 2094 2131
rect 2274 2128 2334 2131
rect 2386 2128 2414 2131
rect 2434 2128 2462 2131
rect 2546 2128 2558 2131
rect 2634 2128 2790 2131
rect 3098 2128 3169 2131
rect 3210 2128 3278 2131
rect 3418 2128 3446 2131
rect 3466 2128 3582 2131
rect 3694 2131 3697 2138
rect 3694 2128 3758 2131
rect 3814 2131 3817 2138
rect 3778 2128 3817 2131
rect 3842 2128 3854 2131
rect 3890 2128 3926 2131
rect 4066 2128 4078 2131
rect 4090 2128 4094 2131
rect 4138 2128 4166 2131
rect 4226 2128 4278 2131
rect 4330 2128 4382 2131
rect 1614 2122 1617 2128
rect 2806 2122 2809 2128
rect 50 2118 206 2121
rect 210 2118 294 2121
rect 298 2118 494 2121
rect 498 2118 646 2121
rect 658 2118 974 2121
rect 1146 2118 1174 2121
rect 1178 2118 1606 2121
rect 1706 2118 1742 2121
rect 1810 2118 2126 2121
rect 2130 2118 2542 2121
rect 2562 2118 2654 2121
rect 2678 2118 2686 2121
rect 2690 2118 2710 2121
rect 2910 2121 2913 2128
rect 3166 2121 3169 2128
rect 3326 2121 3329 2128
rect 2910 2118 3161 2121
rect 3166 2118 3329 2121
rect 3362 2118 3390 2121
rect 3394 2118 3566 2121
rect 3614 2121 3617 2128
rect 3614 2118 3734 2121
rect 3822 2121 3825 2128
rect 3822 2118 4126 2121
rect 4250 2118 4302 2121
rect 418 2108 518 2111
rect 546 2108 582 2111
rect 586 2108 614 2111
rect 658 2108 686 2111
rect 810 2108 886 2111
rect 1042 2108 1062 2111
rect 1082 2108 1118 2111
rect 1298 2108 1406 2111
rect 1442 2108 1486 2111
rect 1546 2108 1838 2111
rect 1842 2108 1910 2111
rect 2162 2108 2230 2111
rect 2266 2108 2326 2111
rect 2330 2108 2358 2111
rect 2410 2108 2438 2111
rect 2442 2108 2598 2111
rect 2602 2108 2742 2111
rect 2754 2108 2838 2111
rect 2866 2108 2894 2111
rect 3158 2111 3161 2118
rect 3158 2108 3214 2111
rect 3314 2108 3358 2111
rect 3386 2108 3438 2111
rect 3442 2108 3502 2111
rect 3530 2108 3638 2111
rect 3642 2108 3958 2111
rect 4018 2108 4270 2111
rect 896 2103 898 2107
rect 902 2103 905 2107
rect 910 2103 912 2107
rect 1534 2102 1537 2108
rect 1928 2103 1930 2107
rect 1934 2103 1937 2107
rect 1942 2103 1944 2107
rect 2952 2103 2954 2107
rect 2958 2103 2961 2107
rect 2966 2103 2968 2107
rect 3976 2103 3978 2107
rect 3982 2103 3985 2107
rect 3990 2103 3992 2107
rect 186 2098 686 2101
rect 1050 2098 1054 2101
rect 1066 2098 1198 2101
rect 1234 2098 1494 2101
rect 1498 2098 1518 2101
rect 1698 2098 1710 2101
rect 1762 2098 1886 2101
rect 1954 2098 1974 2101
rect 1994 2098 2022 2101
rect 2026 2098 2062 2101
rect 2066 2098 2150 2101
rect 2218 2098 2286 2101
rect 2322 2098 2342 2101
rect 2386 2098 2398 2101
rect 2402 2098 2470 2101
rect 2530 2098 2638 2101
rect 2650 2098 2862 2101
rect 2866 2098 2902 2101
rect 3138 2098 3206 2101
rect 3222 2098 3310 2101
rect 3338 2098 3462 2101
rect 3714 2098 3806 2101
rect 3810 2098 3878 2101
rect 4066 2098 4078 2101
rect 4082 2098 4150 2101
rect 4170 2098 4198 2101
rect 4202 2098 4294 2101
rect 4362 2098 4374 2101
rect 170 2088 334 2091
rect 450 2088 470 2091
rect 802 2088 862 2091
rect 866 2088 982 2091
rect 1002 2088 1006 2091
rect 1010 2088 1062 2091
rect 1138 2088 1206 2091
rect 1210 2088 1601 2091
rect 166 2082 169 2088
rect 646 2082 649 2088
rect 290 2078 422 2081
rect 434 2078 606 2081
rect 726 2081 729 2088
rect 1598 2082 1601 2088
rect 1842 2088 2086 2091
rect 2114 2088 2246 2091
rect 2618 2088 2622 2091
rect 2706 2088 2710 2091
rect 2738 2088 2862 2091
rect 2890 2088 2910 2091
rect 3170 2088 3174 2091
rect 3178 2088 3190 2091
rect 3222 2091 3225 2098
rect 3202 2088 3225 2091
rect 3258 2088 3265 2091
rect 3274 2088 3302 2091
rect 3310 2091 3313 2098
rect 3310 2088 3382 2091
rect 3498 2088 3542 2091
rect 3714 2088 3718 2091
rect 3730 2088 3822 2091
rect 3938 2088 4030 2091
rect 4070 2088 4190 2091
rect 1710 2082 1713 2088
rect 726 2078 934 2081
rect 946 2078 950 2081
rect 970 2078 1078 2081
rect 1346 2078 1385 2081
rect 34 2068 62 2071
rect 66 2068 78 2071
rect 474 2068 502 2071
rect 506 2068 654 2071
rect 786 2068 790 2071
rect 802 2068 854 2071
rect 862 2068 889 2071
rect 922 2068 990 2071
rect 1182 2071 1185 2078
rect 1270 2071 1273 2078
rect 994 2068 1049 2071
rect 1182 2068 1273 2071
rect 1382 2072 1385 2078
rect 1530 2078 1566 2081
rect 1722 2078 1878 2081
rect 1882 2078 2302 2081
rect 2338 2078 2374 2081
rect 2378 2078 2382 2081
rect 2418 2078 2502 2081
rect 2554 2078 2774 2081
rect 2794 2078 2798 2081
rect 2826 2078 2830 2081
rect 2870 2081 2873 2088
rect 2842 2078 2873 2081
rect 2930 2078 3014 2081
rect 3106 2078 3110 2081
rect 3186 2078 3214 2081
rect 3230 2081 3233 2088
rect 3246 2082 3249 2088
rect 3574 2082 3577 2088
rect 3230 2078 3238 2081
rect 3258 2078 3278 2081
rect 3282 2078 3406 2081
rect 3426 2078 3454 2081
rect 3474 2078 3518 2081
rect 3830 2081 3833 2088
rect 3770 2078 3833 2081
rect 4062 2081 4065 2088
rect 3858 2078 4065 2081
rect 4070 2082 4073 2088
rect 4114 2078 4118 2081
rect 4170 2078 4174 2081
rect 4178 2078 4222 2081
rect 4258 2078 4262 2081
rect 4330 2078 4334 2081
rect 1406 2072 1409 2078
rect 4366 2072 4369 2078
rect 1474 2068 1614 2071
rect 1618 2068 1694 2071
rect 1874 2068 1886 2071
rect 1906 2068 1974 2071
rect 2042 2068 2078 2071
rect 2122 2068 2126 2071
rect 2302 2068 2422 2071
rect 2426 2068 2433 2071
rect 2442 2068 2446 2071
rect 2514 2068 2550 2071
rect 2554 2068 2686 2071
rect 2706 2068 2718 2071
rect 2762 2068 3190 2071
rect 3202 2068 3230 2071
rect 3234 2068 3326 2071
rect 3338 2068 3342 2071
rect 3410 2068 3510 2071
rect 3530 2068 3561 2071
rect 3618 2068 3622 2071
rect 3642 2068 3646 2071
rect 3682 2068 3790 2071
rect 3890 2068 3918 2071
rect 3922 2068 3950 2071
rect 3962 2068 3998 2071
rect 4002 2068 4006 2071
rect 4026 2068 4030 2071
rect 4050 2068 4054 2071
rect 4082 2068 4102 2071
rect 4162 2068 4206 2071
rect 4250 2068 4318 2071
rect 4330 2068 4334 2071
rect 242 2058 246 2061
rect 250 2058 262 2061
rect 322 2058 478 2061
rect 514 2058 526 2061
rect 530 2058 534 2061
rect 594 2058 622 2061
rect 754 2058 758 2061
rect 862 2061 865 2068
rect 818 2058 865 2061
rect 886 2061 889 2068
rect 1046 2062 1049 2068
rect 1726 2062 1729 2068
rect 2158 2062 2161 2068
rect 2302 2062 2305 2068
rect 886 2058 950 2061
rect 954 2058 961 2061
rect 986 2058 1014 2061
rect 1074 2058 1078 2061
rect 1106 2058 1190 2061
rect 1194 2058 1214 2061
rect 1274 2058 1286 2061
rect 1466 2058 1502 2061
rect 1578 2058 1590 2061
rect 1594 2058 1638 2061
rect 1850 2058 1894 2061
rect 1898 2058 2070 2061
rect 2074 2058 2086 2061
rect 2090 2058 2110 2061
rect 2354 2058 2366 2061
rect 2410 2058 2414 2061
rect 2418 2058 2494 2061
rect 2498 2058 2510 2061
rect 2514 2058 2710 2061
rect 2714 2058 2846 2061
rect 2898 2058 2918 2061
rect 3002 2058 3198 2061
rect 3210 2058 3310 2061
rect 3374 2061 3377 2068
rect 3330 2058 3377 2061
rect 3458 2058 3550 2061
rect 3558 2061 3561 2068
rect 3846 2062 3849 2068
rect 3558 2058 3638 2061
rect 3642 2058 3702 2061
rect 3722 2058 3750 2061
rect 3890 2058 3894 2061
rect 3946 2058 4105 2061
rect 4114 2058 4142 2061
rect 4146 2058 4358 2061
rect 4362 2058 4366 2061
rect 782 2052 785 2058
rect 878 2052 881 2058
rect 3814 2052 3817 2058
rect -26 2051 -22 2052
rect -26 2048 6 2051
rect 58 2048 86 2051
rect 522 2048 526 2051
rect 622 2048 630 2051
rect 634 2048 662 2051
rect 666 2048 678 2051
rect 722 2048 766 2051
rect 770 2048 774 2051
rect 882 2048 1126 2051
rect 1162 2048 1166 2051
rect 1194 2048 1198 2051
rect 1362 2048 1566 2051
rect 1826 2048 1934 2051
rect 1938 2048 1942 2051
rect 1970 2048 2014 2051
rect 2058 2048 2126 2051
rect 2130 2048 2142 2051
rect 2530 2048 2534 2051
rect 2554 2048 2582 2051
rect 2730 2048 2753 2051
rect 2762 2048 2766 2051
rect 2778 2048 2782 2051
rect 2790 2048 2809 2051
rect 3090 2048 3166 2051
rect 3242 2048 3262 2051
rect 3282 2048 3294 2051
rect 3330 2048 3350 2051
rect 3354 2048 3366 2051
rect 3410 2048 3414 2051
rect 3466 2048 3486 2051
rect 3594 2048 3702 2051
rect 3758 2048 3774 2051
rect 4018 2048 4062 2051
rect 4102 2051 4105 2058
rect 4102 2048 4206 2051
rect 4306 2048 4337 2051
rect 2750 2042 2753 2048
rect 2790 2042 2793 2048
rect 2806 2042 2809 2048
rect 3710 2042 3713 2048
rect 3758 2042 3761 2048
rect 4334 2042 4337 2048
rect 490 2038 742 2041
rect 754 2038 806 2041
rect 810 2038 822 2041
rect 890 2038 982 2041
rect 986 2038 1110 2041
rect 1126 2038 1142 2041
rect 1178 2038 1382 2041
rect 1386 2038 1494 2041
rect 1522 2038 1782 2041
rect 1866 2038 1870 2041
rect 1882 2038 1998 2041
rect 2010 2038 2662 2041
rect 2826 2038 2910 2041
rect 3138 2038 3246 2041
rect 3346 2038 3518 2041
rect 3578 2038 3606 2041
rect 3610 2038 3630 2041
rect 3802 2038 3910 2041
rect 3914 2038 4046 2041
rect 4050 2038 4118 2041
rect 4274 2038 4302 2041
rect 1126 2032 1129 2038
rect 682 2028 774 2031
rect 938 2028 990 2031
rect 994 2028 1014 2031
rect 1034 2028 1086 2031
rect 1146 2028 1398 2031
rect 1442 2028 1902 2031
rect 1906 2028 2478 2031
rect 2482 2028 2534 2031
rect 2538 2028 2574 2031
rect 2682 2028 2798 2031
rect 2802 2028 3126 2031
rect 3210 2028 3230 2031
rect 3342 2031 3345 2038
rect 3234 2028 3345 2031
rect 3526 2031 3529 2038
rect 4150 2032 4153 2038
rect 3526 2028 3782 2031
rect 4018 2028 4094 2031
rect 806 2021 809 2028
rect 690 2018 809 2021
rect 818 2018 942 2021
rect 946 2018 1118 2021
rect 1154 2018 1230 2021
rect 1234 2018 1350 2021
rect 1398 2021 1401 2028
rect 1398 2018 2734 2021
rect 2746 2018 2750 2021
rect 2770 2018 3086 2021
rect 3098 2018 3390 2021
rect 3394 2018 3598 2021
rect 3602 2018 3854 2021
rect -26 2011 -22 2012
rect -26 2008 6 2011
rect 634 2008 638 2011
rect 662 2008 942 2011
rect 946 2008 1006 2011
rect 1034 2008 1102 2011
rect 1130 2008 1158 2011
rect 1466 2008 1646 2011
rect 1834 2008 1838 2011
rect 1850 2008 1862 2011
rect 1866 2008 1878 2011
rect 1890 2008 1894 2011
rect 2034 2008 2038 2011
rect 2050 2008 2206 2011
rect 2210 2008 2398 2011
rect 2618 2008 2638 2011
rect 2650 2008 2822 2011
rect 2826 2008 2926 2011
rect 2930 2008 3054 2011
rect 3058 2008 3462 2011
rect 3586 2008 3654 2011
rect 3850 2008 3942 2011
rect 3946 2008 3950 2011
rect 4138 2008 4238 2011
rect 392 2003 394 2007
rect 398 2003 401 2007
rect 406 2003 408 2007
rect 662 2002 665 2008
rect 1416 2003 1418 2007
rect 1422 2003 1425 2007
rect 1430 2003 1432 2007
rect 2440 2003 2442 2007
rect 2446 2003 2449 2007
rect 2454 2003 2456 2007
rect 3472 2003 3474 2007
rect 3478 2003 3481 2007
rect 3486 2003 3488 2007
rect 10 1998 142 2001
rect 626 1998 662 2001
rect 674 1998 694 2001
rect 706 1998 766 2001
rect 778 1998 830 2001
rect 866 1998 977 2001
rect 1042 1998 1054 2001
rect 1162 1998 1390 2001
rect 1554 1998 1558 2001
rect 1602 1998 1614 2001
rect 1622 1998 1966 2001
rect 2074 1998 2174 2001
rect 2186 1998 2198 2001
rect 2634 1998 2846 2001
rect 2850 1998 2934 2001
rect 3186 1998 3286 2001
rect 3298 1998 3310 2001
rect 3362 1998 3430 2001
rect 3594 1998 4230 2001
rect -26 1991 -22 1992
rect -26 1988 38 1991
rect 74 1988 702 1991
rect 706 1988 774 1991
rect 818 1988 822 1991
rect 858 1988 878 1991
rect 882 1988 934 1991
rect 974 1991 977 1998
rect 974 1988 1078 1991
rect 1622 1991 1625 1998
rect 1386 1988 1625 1991
rect 1634 1988 1678 1991
rect 1738 1988 1750 1991
rect 1778 1988 1806 1991
rect 1830 1988 1838 1991
rect 1842 1988 1854 1991
rect 1862 1988 1870 1991
rect 1874 1988 1942 1991
rect 1962 1988 2662 1991
rect 2666 1988 2950 1991
rect 3214 1988 3398 1991
rect 3530 1988 3622 1991
rect -26 1978 126 1981
rect 226 1978 446 1981
rect 690 1978 742 1981
rect 778 1978 870 1981
rect 986 1978 990 1981
rect 1002 1978 1102 1981
rect 1262 1981 1265 1988
rect 1318 1982 1321 1988
rect 3214 1982 3217 1988
rect 1186 1978 1265 1981
rect 1346 1978 1454 1981
rect 1474 1978 1966 1981
rect 1978 1978 2158 1981
rect 2666 1978 3006 1981
rect 3098 1978 3214 1981
rect 3278 1978 3286 1981
rect 3290 1978 3414 1981
rect 3650 1978 3758 1981
rect -26 1972 -23 1978
rect -26 1968 -22 1972
rect 82 1968 230 1971
rect 638 1971 641 1978
rect 354 1968 641 1971
rect 658 1968 670 1971
rect 690 1968 694 1971
rect 714 1968 718 1971
rect 730 1968 758 1971
rect 762 1968 822 1971
rect 926 1971 929 1978
rect 850 1968 929 1971
rect 954 1968 1014 1971
rect 1018 1968 1070 1971
rect 1258 1968 1262 1971
rect 1302 1971 1305 1978
rect 1282 1968 1305 1971
rect 1314 1968 1542 1971
rect 1610 1968 1718 1971
rect 1778 1968 1798 1971
rect 2074 1968 2558 1971
rect 2562 1968 2574 1971
rect 2582 1971 2585 1978
rect 4166 1972 4169 1978
rect 2582 1968 2622 1971
rect 2626 1968 2790 1971
rect 2946 1968 3062 1971
rect 3066 1968 3094 1971
rect 3186 1968 3342 1971
rect 3386 1968 3430 1971
rect 3514 1968 3622 1971
rect 3770 1968 3918 1971
rect 4138 1968 4142 1971
rect 4214 1971 4217 1978
rect 4294 1972 4297 1978
rect 4214 1968 4230 1971
rect 62 1961 65 1968
rect 26 1958 65 1961
rect 74 1958 102 1961
rect 138 1958 182 1961
rect 238 1961 241 1968
rect 238 1958 638 1961
rect 642 1958 726 1961
rect 786 1958 998 1961
rect 1002 1958 1022 1961
rect 1138 1958 1142 1961
rect 1162 1958 1166 1961
rect 1266 1958 1374 1961
rect 1378 1958 1438 1961
rect 1982 1961 1985 1968
rect 1578 1958 1985 1961
rect 2002 1958 2118 1961
rect 2482 1958 2510 1961
rect 2634 1958 2638 1961
rect 2818 1958 3070 1961
rect 3090 1958 3110 1961
rect 3170 1958 3206 1961
rect 3218 1958 3406 1961
rect 3426 1958 3542 1961
rect 3546 1958 3553 1961
rect 3562 1958 3606 1961
rect 3682 1958 3702 1961
rect 3954 1958 4006 1961
rect 4154 1958 4254 1961
rect 4274 1958 4310 1961
rect 206 1952 209 1958
rect 2590 1952 2593 1958
rect 3606 1952 3609 1958
rect 4094 1952 4097 1958
rect 4342 1952 4345 1958
rect -26 1951 -22 1952
rect -26 1948 6 1951
rect 58 1948 62 1951
rect 74 1948 102 1951
rect 106 1948 174 1951
rect 546 1948 678 1951
rect 710 1948 718 1951
rect 794 1948 798 1951
rect 810 1948 814 1951
rect 842 1948 862 1951
rect 874 1948 966 1951
rect 970 1948 1030 1951
rect 1034 1948 1054 1951
rect 1074 1948 1166 1951
rect 1218 1948 1278 1951
rect 1330 1948 1366 1951
rect 1386 1948 1574 1951
rect 1722 1948 1742 1951
rect 1754 1948 1785 1951
rect 1802 1948 1926 1951
rect 1938 1948 2014 1951
rect 2170 1948 2174 1951
rect 2282 1948 2366 1951
rect 2506 1948 2518 1951
rect 2770 1948 2782 1951
rect 2826 1948 2886 1951
rect 3002 1948 3046 1951
rect 3130 1948 3137 1951
rect 3146 1948 3150 1951
rect 3202 1948 3222 1951
rect 3346 1948 3350 1951
rect 3442 1948 3446 1951
rect 3562 1948 3590 1951
rect 3722 1948 3734 1951
rect 3962 1948 4014 1951
rect 4082 1948 4094 1951
rect 4130 1948 4142 1951
rect 4210 1948 4294 1951
rect 174 1942 177 1948
rect 162 1938 166 1941
rect 194 1938 222 1941
rect 254 1941 257 1948
rect 710 1942 713 1948
rect 1782 1942 1785 1948
rect 2038 1942 2041 1948
rect 234 1938 257 1941
rect 458 1938 614 1941
rect 642 1938 654 1941
rect 690 1938 702 1941
rect 746 1938 910 1941
rect 930 1938 982 1941
rect 994 1938 998 1941
rect 1026 1938 1030 1941
rect 1090 1938 1134 1941
rect 1146 1938 1150 1941
rect 1162 1938 1166 1941
rect 1242 1938 1246 1941
rect 1274 1938 1278 1941
rect 1282 1938 1350 1941
rect 1362 1938 1366 1941
rect 1442 1938 1446 1941
rect 1738 1938 1758 1941
rect 1906 1938 1910 1941
rect 1922 1938 1990 1941
rect 2234 1938 2326 1941
rect 2382 1941 2385 1948
rect 2486 1941 2489 1948
rect 2942 1942 2945 1948
rect 2382 1938 2489 1941
rect 2526 1938 2598 1941
rect 2666 1938 2726 1941
rect 2730 1938 2902 1941
rect 2978 1938 3022 1941
rect 3026 1938 3086 1941
rect 3122 1938 3174 1941
rect 3178 1938 3182 1941
rect 3258 1938 3262 1941
rect 3274 1938 3310 1941
rect 3314 1938 3318 1941
rect 3322 1938 3358 1941
rect 3410 1938 3462 1941
rect 3514 1938 3526 1941
rect 3534 1941 3537 1948
rect 3534 1938 3614 1941
rect 3622 1941 3625 1948
rect 3622 1938 3670 1941
rect 3698 1938 3718 1941
rect 3722 1938 3742 1941
rect 3862 1941 3865 1948
rect 4038 1942 4041 1948
rect 3786 1938 3865 1941
rect 3938 1938 3966 1941
rect 4042 1938 4070 1941
rect 4082 1938 4086 1941
rect 4114 1938 4166 1941
rect 4178 1938 4182 1941
rect 4202 1938 4214 1941
rect 4258 1938 4278 1941
rect 4330 1938 4366 1941
rect 334 1932 337 1938
rect 90 1928 166 1931
rect 170 1928 198 1931
rect 714 1928 1198 1931
rect 1202 1928 1302 1931
rect 1330 1928 1342 1931
rect 1390 1931 1393 1938
rect 1354 1928 1393 1931
rect 1442 1928 1462 1931
rect 1482 1928 1486 1931
rect 1590 1931 1593 1938
rect 1806 1932 1809 1938
rect 2014 1932 2017 1938
rect 2166 1932 2169 1938
rect 1586 1928 1593 1931
rect 1618 1928 1678 1931
rect 2226 1928 2246 1931
rect 2250 1928 2270 1931
rect 2282 1928 2358 1931
rect 2366 1931 2369 1938
rect 2362 1928 2369 1931
rect 2526 1931 2529 1938
rect 2434 1928 2529 1931
rect 2538 1928 2670 1931
rect 2674 1928 2686 1931
rect 2750 1928 2806 1931
rect 2810 1928 2870 1931
rect 3054 1928 3062 1931
rect 3066 1928 3078 1931
rect 3086 1928 3094 1931
rect 3098 1928 3150 1931
rect 3162 1928 3206 1931
rect 3258 1928 3278 1931
rect 3290 1928 3318 1931
rect 3322 1928 3398 1931
rect 3546 1928 3590 1931
rect 3602 1928 3630 1931
rect 3634 1928 3646 1931
rect 3650 1928 3798 1931
rect 3850 1928 4014 1931
rect 4162 1928 4182 1931
rect 4226 1928 4262 1931
rect 4306 1928 4350 1931
rect 4354 1928 4390 1931
rect 526 1922 529 1928
rect 2750 1922 2753 1928
rect 194 1918 262 1921
rect 770 1918 782 1921
rect 786 1918 793 1921
rect 826 1918 1238 1921
rect 1242 1918 1662 1921
rect 1670 1918 1742 1921
rect 1746 1918 1758 1921
rect 1770 1918 1798 1921
rect 2002 1918 2030 1921
rect 2186 1918 2273 1921
rect 2282 1918 2454 1921
rect 2466 1918 2566 1921
rect 2610 1918 2750 1921
rect 3066 1918 3102 1921
rect 3130 1918 3182 1921
rect 3282 1918 3438 1921
rect 3578 1918 3622 1921
rect 3682 1918 3726 1921
rect 3754 1918 3894 1921
rect 4086 1921 4089 1928
rect 3898 1918 4089 1921
rect 4290 1918 4302 1921
rect 4346 1918 4358 1921
rect 1670 1912 1673 1918
rect 370 1908 526 1911
rect 602 1908 630 1911
rect 634 1908 886 1911
rect 978 1908 1102 1911
rect 1114 1908 1118 1911
rect 1146 1908 1222 1911
rect 1314 1908 1382 1911
rect 1394 1908 1406 1911
rect 1450 1908 1478 1911
rect 1570 1908 1598 1911
rect 1610 1908 1654 1911
rect 1706 1908 1814 1911
rect 1850 1908 1854 1911
rect 1858 1908 1918 1911
rect 2058 1908 2078 1911
rect 2138 1908 2262 1911
rect 2270 1911 2273 1918
rect 2270 1908 2294 1911
rect 2362 1908 2382 1911
rect 2418 1908 2430 1911
rect 2434 1908 2502 1911
rect 2566 1911 2569 1918
rect 2566 1908 2726 1911
rect 2730 1908 2814 1911
rect 3170 1908 3350 1911
rect 3458 1908 3510 1911
rect 3514 1908 3582 1911
rect 3706 1908 3878 1911
rect 3906 1908 3910 1911
rect 4066 1908 4102 1911
rect 4290 1908 4310 1911
rect 896 1903 898 1907
rect 902 1903 905 1907
rect 910 1903 912 1907
rect 1928 1903 1930 1907
rect 1934 1903 1937 1907
rect 1942 1903 1944 1907
rect 2952 1903 2954 1907
rect 2958 1903 2961 1907
rect 2966 1903 2968 1907
rect 3976 1903 3978 1907
rect 3982 1903 3985 1907
rect 3990 1903 3992 1907
rect 66 1898 206 1901
rect 402 1898 430 1901
rect 538 1898 806 1901
rect 874 1898 886 1901
rect 978 1898 1462 1901
rect 1482 1898 1510 1901
rect 1618 1898 1630 1901
rect 1666 1898 1774 1901
rect 1898 1898 1902 1901
rect 2026 1898 2126 1901
rect 2130 1898 2430 1901
rect 2442 1898 2654 1901
rect 2778 1898 2790 1901
rect 2986 1898 3118 1901
rect 3146 1898 3174 1901
rect 3226 1898 3294 1901
rect 3298 1898 3334 1901
rect 3450 1898 3494 1901
rect 3522 1898 3646 1901
rect 3650 1898 3934 1901
rect 4226 1898 4246 1901
rect 114 1888 286 1891
rect 290 1888 294 1891
rect 426 1888 1014 1891
rect 1018 1888 1158 1891
rect 1162 1888 1366 1891
rect 1570 1888 1574 1891
rect 1618 1888 1646 1891
rect 1914 1888 1918 1891
rect 1922 1888 2118 1891
rect 2186 1888 2233 1891
rect 2306 1888 2382 1891
rect 2682 1888 2718 1891
rect 3114 1888 3126 1891
rect 3130 1888 3137 1891
rect 3162 1888 3214 1891
rect 3218 1888 3518 1891
rect 3530 1888 3542 1891
rect 3702 1888 3710 1891
rect 3738 1888 3742 1891
rect 3746 1888 3806 1891
rect 3810 1888 3886 1891
rect 3914 1888 4006 1891
rect 4154 1888 4281 1891
rect 4298 1888 4310 1891
rect 1470 1882 1473 1888
rect 1766 1882 1769 1888
rect 58 1878 86 1881
rect 90 1878 102 1881
rect 658 1878 726 1881
rect 778 1878 854 1881
rect 866 1878 902 1881
rect 1034 1878 1038 1881
rect 1114 1878 1126 1881
rect 1138 1878 1214 1881
rect 1258 1878 1294 1881
rect 1322 1878 1334 1881
rect 1410 1878 1454 1881
rect 1530 1878 1630 1881
rect 1634 1878 1686 1881
rect 1870 1881 1873 1888
rect 2230 1882 2233 1888
rect 1870 1878 1878 1881
rect 1922 1878 2006 1881
rect 2090 1878 2094 1881
rect 2130 1878 2214 1881
rect 2398 1881 2401 1888
rect 2398 1878 2430 1881
rect 2434 1878 2478 1881
rect 2590 1881 2593 1888
rect 4278 1882 4281 1888
rect 2522 1878 2593 1881
rect 2610 1878 2809 1881
rect 2930 1878 2950 1881
rect 2954 1878 2974 1881
rect 3002 1878 3417 1881
rect -26 1871 -22 1872
rect 30 1871 33 1878
rect -26 1868 33 1871
rect 190 1872 193 1878
rect 382 1872 385 1878
rect 534 1872 537 1878
rect 550 1872 553 1878
rect 774 1872 777 1878
rect 1006 1872 1009 1878
rect 1510 1872 1513 1878
rect 822 1868 830 1871
rect 834 1868 838 1871
rect 866 1868 870 1871
rect 890 1868 958 1871
rect 1010 1868 1174 1871
rect 1178 1868 1326 1871
rect 1330 1868 1494 1871
rect 1518 1868 1702 1871
rect 1954 1868 2022 1871
rect 2054 1871 2057 1878
rect 2054 1868 2198 1871
rect 2262 1870 2334 1871
rect 34 1858 70 1861
rect 442 1858 478 1861
rect 710 1861 713 1868
rect 706 1858 713 1861
rect 730 1858 734 1861
rect 778 1858 782 1861
rect 802 1858 822 1861
rect 850 1858 862 1861
rect 882 1858 918 1861
rect 970 1858 982 1861
rect 1010 1858 1038 1861
rect 1042 1858 1054 1861
rect 1074 1858 1078 1861
rect 1098 1858 1110 1861
rect 1146 1858 1206 1861
rect 1226 1858 1270 1861
rect 1282 1858 1286 1861
rect 1298 1858 1302 1861
rect 1362 1858 1462 1861
rect 1518 1861 1521 1868
rect 1726 1862 1729 1868
rect 2266 1868 2334 1870
rect 2514 1868 2678 1871
rect 2806 1871 2809 1878
rect 3414 1872 3417 1878
rect 3498 1878 3542 1881
rect 3562 1878 3702 1881
rect 3706 1878 3742 1881
rect 3770 1878 3790 1881
rect 3802 1878 3814 1881
rect 3818 1878 3862 1881
rect 3866 1878 3958 1881
rect 4074 1878 4078 1881
rect 4170 1878 4230 1881
rect 2794 1868 2801 1871
rect 2806 1868 3086 1871
rect 3090 1868 3097 1871
rect 3106 1868 3182 1871
rect 3202 1868 3238 1871
rect 3430 1871 3433 1878
rect 4142 1872 4145 1878
rect 3430 1868 3526 1871
rect 3538 1868 3550 1871
rect 3602 1868 3726 1871
rect 3730 1868 3774 1871
rect 3802 1868 3942 1871
rect 4002 1868 4022 1871
rect 4194 1868 4318 1871
rect 4322 1868 4326 1871
rect 4338 1868 4366 1871
rect 2366 1862 2369 1868
rect 1466 1858 1521 1861
rect 1554 1858 1566 1861
rect 1650 1858 1673 1861
rect 1698 1858 1705 1861
rect 1746 1858 1750 1861
rect 2010 1858 2030 1861
rect 2074 1858 2089 1861
rect 1534 1852 1537 1858
rect 1670 1852 1673 1858
rect 1702 1852 1705 1858
rect 2054 1852 2057 1858
rect 2086 1852 2089 1858
rect 2098 1858 2142 1861
rect 2146 1858 2246 1861
rect 2298 1858 2318 1861
rect 2406 1861 2409 1868
rect 2798 1862 2801 1868
rect 2386 1858 2409 1861
rect 2474 1858 2478 1861
rect 2506 1858 2542 1861
rect 2666 1858 2694 1861
rect 2714 1858 2734 1861
rect 2818 1858 2878 1861
rect 2882 1858 2942 1861
rect 2946 1858 2974 1861
rect 3082 1858 3150 1861
rect 3178 1858 3206 1861
rect 3210 1858 3246 1861
rect 3330 1858 3510 1861
rect 3562 1858 3606 1861
rect 3626 1858 3694 1861
rect 3698 1858 3734 1861
rect 3754 1858 3758 1861
rect 3794 1858 3822 1861
rect 3922 1858 3942 1861
rect 3978 1858 3990 1861
rect 4082 1858 4086 1861
rect 4106 1858 4110 1861
rect 4130 1858 4150 1861
rect 4258 1858 4310 1861
rect 4342 1858 4358 1861
rect 2094 1852 2097 1858
rect -26 1851 -22 1852
rect -26 1848 6 1851
rect 58 1848 86 1851
rect 178 1848 550 1851
rect 702 1848 758 1851
rect 898 1848 1462 1851
rect 1466 1848 1470 1851
rect 1642 1848 1654 1851
rect 1658 1848 1662 1851
rect 1726 1848 1854 1851
rect 2106 1848 2166 1851
rect 2226 1848 2246 1851
rect 2258 1848 2342 1851
rect 2346 1848 2462 1851
rect 2690 1848 2718 1851
rect 2806 1851 2809 1858
rect 4238 1852 4241 1858
rect 4342 1852 4345 1858
rect 2722 1848 2777 1851
rect 2806 1848 3078 1851
rect 3090 1848 3190 1851
rect 3602 1848 3630 1851
rect 3658 1848 3678 1851
rect 3738 1848 3774 1851
rect 3834 1848 3894 1851
rect 4002 1848 4198 1851
rect 4250 1848 4326 1851
rect 702 1842 705 1848
rect 282 1838 654 1841
rect 782 1841 785 1848
rect 746 1838 785 1841
rect 794 1838 1134 1841
rect 1226 1838 1254 1841
rect 1370 1838 1374 1841
rect 1418 1838 1422 1841
rect 1450 1838 1454 1841
rect 1482 1838 1494 1841
rect 1498 1838 1550 1841
rect 1726 1841 1729 1848
rect 2774 1842 2777 1848
rect 1642 1838 1729 1841
rect 1738 1838 2406 1841
rect 2410 1838 2534 1841
rect 2538 1838 2646 1841
rect 2658 1838 2694 1841
rect 2698 1838 2742 1841
rect 2778 1838 2798 1841
rect 3018 1838 3310 1841
rect 3314 1838 3326 1841
rect 3674 1838 3774 1841
rect 3778 1838 3830 1841
rect 3834 1838 3918 1841
rect 3930 1838 3950 1841
rect 4166 1838 4174 1841
rect 4202 1838 4246 1841
rect 4166 1832 4169 1838
rect 82 1828 462 1831
rect 778 1828 830 1831
rect 914 1828 918 1831
rect 978 1828 998 1831
rect 1034 1828 1105 1831
rect 1170 1828 1262 1831
rect 1338 1828 1342 1831
rect 1362 1828 1382 1831
rect 1394 1828 1582 1831
rect 1586 1828 1630 1831
rect 1634 1828 1694 1831
rect 1962 1828 3694 1831
rect 3706 1828 3718 1831
rect 3722 1828 4062 1831
rect 4274 1828 4294 1831
rect 4298 1828 4382 1831
rect 474 1818 798 1821
rect 802 1818 806 1821
rect 818 1818 830 1821
rect 834 1818 870 1821
rect 974 1821 977 1828
rect 1102 1822 1105 1828
rect 874 1818 977 1821
rect 1066 1818 1078 1821
rect 1138 1818 1318 1821
rect 1350 1821 1353 1828
rect 1346 1818 1353 1821
rect 1378 1818 1854 1821
rect 1994 1818 2070 1821
rect 2082 1818 2326 1821
rect 2330 1818 2390 1821
rect 2506 1818 2510 1821
rect 2530 1818 2662 1821
rect 2666 1818 2750 1821
rect 2762 1818 2846 1821
rect 3030 1818 3038 1821
rect 3042 1818 3054 1821
rect 3122 1818 3142 1821
rect 3258 1818 3374 1821
rect 3410 1818 3534 1821
rect 3666 1818 3710 1821
rect 3714 1818 3742 1821
rect 3754 1818 3870 1821
rect 3878 1818 4062 1821
rect 690 1808 742 1811
rect 802 1808 958 1811
rect 962 1808 1222 1811
rect 1234 1808 1406 1811
rect 1442 1808 1486 1811
rect 1634 1808 1758 1811
rect 1898 1808 2070 1811
rect 2106 1808 2278 1811
rect 2658 1808 3238 1811
rect 3242 1808 3278 1811
rect 3362 1808 3382 1811
rect 3530 1808 3750 1811
rect 3878 1811 3881 1818
rect 3754 1808 3881 1811
rect 392 1803 394 1807
rect 398 1803 401 1807
rect 406 1803 408 1807
rect 1416 1803 1418 1807
rect 1422 1803 1425 1807
rect 1430 1803 1432 1807
rect 2440 1803 2442 1807
rect 2446 1803 2449 1807
rect 2454 1803 2456 1807
rect 3472 1803 3474 1807
rect 3478 1803 3481 1807
rect 3486 1803 3488 1807
rect 506 1798 1270 1801
rect 1354 1798 1374 1801
rect 1594 1798 1654 1801
rect 1690 1798 1790 1801
rect 1818 1798 2078 1801
rect 2170 1798 2174 1801
rect 2178 1798 2406 1801
rect 2466 1798 2878 1801
rect 3050 1798 3062 1801
rect 3066 1798 3190 1801
rect 3554 1798 3598 1801
rect 3762 1798 3894 1801
rect 3930 1798 4022 1801
rect 4042 1798 4046 1801
rect 4066 1798 4126 1801
rect 4130 1798 4150 1801
rect 4154 1798 4158 1801
rect -26 1791 -22 1792
rect -26 1788 6 1791
rect 250 1788 262 1791
rect 706 1788 1150 1791
rect 1186 1788 1206 1791
rect 1222 1788 1230 1791
rect 1234 1788 1262 1791
rect 1274 1788 2518 1791
rect 2522 1788 2606 1791
rect 2650 1788 3646 1791
rect 3746 1788 3761 1791
rect 4042 1788 4086 1791
rect 4094 1788 4102 1791
rect 4106 1788 4185 1791
rect 4194 1788 4206 1791
rect 3758 1782 3761 1788
rect 658 1778 846 1781
rect 858 1778 1230 1781
rect 1290 1778 1326 1781
rect 1330 1778 1537 1781
rect 1554 1778 1614 1781
rect 1658 1778 1745 1781
rect -26 1771 -22 1772
rect 30 1771 33 1778
rect 1534 1772 1537 1778
rect 1742 1772 1745 1778
rect 1982 1778 2054 1781
rect 2066 1778 2110 1781
rect 2186 1778 2190 1781
rect 2322 1778 2878 1781
rect 3218 1778 3270 1781
rect 3282 1778 3374 1781
rect 3426 1778 3662 1781
rect 3730 1778 3734 1781
rect 3954 1778 3966 1781
rect 3970 1778 4126 1781
rect 4130 1778 4166 1781
rect 4182 1781 4185 1788
rect 4182 1778 4278 1781
rect 4298 1778 4358 1781
rect 1774 1772 1777 1778
rect 1982 1772 1985 1778
rect -26 1768 33 1771
rect 338 1768 662 1771
rect 698 1768 734 1771
rect 890 1768 934 1771
rect 938 1768 950 1771
rect 986 1768 1062 1771
rect 1114 1768 1126 1771
rect 1130 1768 1182 1771
rect 1186 1768 1302 1771
rect 1306 1768 1430 1771
rect 1538 1768 1734 1771
rect 1786 1768 1838 1771
rect 1858 1768 1958 1771
rect 2154 1768 2158 1771
rect 2186 1768 2358 1771
rect 2490 1768 2814 1771
rect 2866 1768 3366 1771
rect 3410 1768 3430 1771
rect 3602 1768 3633 1771
rect 3642 1768 3750 1771
rect 3754 1768 3782 1771
rect 4042 1768 4046 1771
rect 4090 1768 4102 1771
rect 4134 1768 4158 1771
rect 1510 1762 1513 1768
rect 26 1758 438 1761
rect 458 1758 790 1761
rect 978 1758 1006 1761
rect 1026 1758 1070 1761
rect 1130 1758 1142 1761
rect 1154 1758 1158 1761
rect 1202 1758 1246 1761
rect 1250 1758 1302 1761
rect 1306 1758 1454 1761
rect 1458 1758 1486 1761
rect 1522 1758 1662 1761
rect 1682 1758 1729 1761
rect 1738 1758 1990 1761
rect 2070 1761 2073 1768
rect 2058 1758 2073 1761
rect 2078 1762 2081 1768
rect 2154 1758 2190 1761
rect 2226 1758 2230 1761
rect 2242 1758 2246 1761
rect 2274 1758 2454 1761
rect 2478 1761 2481 1768
rect 2478 1758 2534 1761
rect 2586 1758 2590 1761
rect 2658 1758 2702 1761
rect 2706 1758 2710 1761
rect 2738 1758 2758 1761
rect 2770 1758 2790 1761
rect 2826 1758 3014 1761
rect 3098 1758 3102 1761
rect 3146 1758 3174 1761
rect 3186 1758 3294 1761
rect 3370 1758 3454 1761
rect 3458 1758 3614 1761
rect 3630 1761 3633 1768
rect 4134 1762 4137 1768
rect 4174 1762 4177 1768
rect 3630 1758 3678 1761
rect 3682 1758 3734 1761
rect 3794 1758 3974 1761
rect 3994 1758 4006 1761
rect 4010 1758 4054 1761
rect 4058 1758 4110 1761
rect 4114 1758 4118 1761
rect 4146 1758 4158 1761
rect 4342 1761 4345 1768
rect 4194 1758 4345 1761
rect 1726 1752 1729 1758
rect -26 1751 -22 1752
rect -26 1748 6 1751
rect 618 1748 654 1751
rect 890 1748 910 1751
rect 930 1748 1270 1751
rect 1298 1748 1326 1751
rect 1346 1748 1374 1751
rect 1386 1748 1414 1751
rect 1490 1748 1494 1751
rect 1498 1748 1606 1751
rect 1626 1748 1662 1751
rect 1674 1748 1689 1751
rect 2046 1751 2049 1758
rect 1786 1748 2049 1751
rect 2058 1748 2062 1751
rect 2154 1748 2310 1751
rect 2314 1748 2462 1751
rect 2466 1748 2630 1751
rect 2634 1748 2822 1751
rect 2906 1748 3086 1751
rect 3122 1748 3126 1751
rect 3170 1748 3190 1751
rect 3250 1748 3278 1751
rect 3294 1748 3326 1751
rect 3354 1748 3462 1751
rect 3594 1748 3654 1751
rect 3658 1748 3670 1751
rect 3770 1748 3774 1751
rect 3946 1748 3958 1751
rect 3962 1748 4126 1751
rect 4130 1748 4134 1751
rect 4182 1751 4185 1758
rect 4390 1752 4393 1758
rect 4138 1748 4214 1751
rect 4250 1748 4254 1751
rect 4370 1748 4390 1751
rect 158 1742 161 1748
rect 1686 1742 1689 1748
rect 754 1738 830 1741
rect 874 1738 942 1741
rect 946 1738 990 1741
rect 994 1738 1038 1741
rect 1050 1738 1118 1741
rect 1178 1738 1198 1741
rect 1218 1738 1246 1741
rect 1362 1738 1550 1741
rect 1554 1738 1638 1741
rect 1714 1738 1974 1741
rect 2002 1738 2070 1741
rect 2162 1738 2166 1741
rect 2186 1738 2190 1741
rect 2202 1738 2214 1741
rect 2250 1738 2254 1741
rect 2354 1738 2358 1741
rect 2374 1738 2558 1741
rect 2586 1738 2606 1741
rect 2610 1738 2750 1741
rect 2770 1738 2798 1741
rect 3122 1738 3150 1741
rect 3230 1741 3233 1748
rect 3294 1742 3297 1748
rect 3726 1742 3729 1748
rect 3186 1738 3233 1741
rect 3242 1738 3270 1741
rect 3338 1738 3398 1741
rect 3434 1738 3510 1741
rect 3514 1738 3558 1741
rect 3770 1738 3774 1741
rect 4098 1738 4102 1741
rect 4146 1738 4190 1741
rect 142 1731 145 1738
rect 142 1728 270 1731
rect 542 1731 545 1738
rect 274 1728 321 1731
rect 542 1728 574 1731
rect 710 1731 713 1738
rect 1982 1732 1985 1738
rect 2102 1732 2105 1738
rect 2374 1732 2377 1738
rect 3614 1732 3617 1738
rect 3702 1732 3705 1738
rect 710 1728 718 1731
rect 786 1728 806 1731
rect 842 1728 902 1731
rect 922 1728 950 1731
rect 970 1728 990 1731
rect 1018 1728 1054 1731
rect 1058 1728 1062 1731
rect 1074 1728 1078 1731
rect 1210 1728 1230 1731
rect 1250 1728 1262 1731
rect 1330 1728 1366 1731
rect 1370 1728 1526 1731
rect 1546 1728 1558 1731
rect 1586 1728 1694 1731
rect 1698 1728 1702 1731
rect 1850 1728 1873 1731
rect 1890 1728 1958 1731
rect 1994 1728 2006 1731
rect 2014 1728 2022 1731
rect 2026 1728 2030 1731
rect 2050 1728 2086 1731
rect 2122 1728 2230 1731
rect 2690 1728 2710 1731
rect 2746 1728 2774 1731
rect 2786 1728 2838 1731
rect 2842 1728 3126 1731
rect 3146 1728 3278 1731
rect 3282 1728 3582 1731
rect 3586 1728 3590 1731
rect 4050 1728 4166 1731
rect 4170 1728 4190 1731
rect 4202 1728 4222 1731
rect 318 1722 321 1728
rect 950 1722 953 1728
rect 1870 1722 1873 1728
rect 474 1718 486 1721
rect 530 1718 542 1721
rect 698 1718 862 1721
rect 930 1718 934 1721
rect 970 1718 1014 1721
rect 1026 1718 1038 1721
rect 1074 1718 1166 1721
rect 1334 1718 1342 1721
rect 1346 1718 1366 1721
rect 1394 1718 1398 1721
rect 1538 1718 1558 1721
rect 1602 1718 1678 1721
rect 1786 1718 1790 1721
rect 1810 1718 1814 1721
rect 1918 1718 2270 1721
rect 2370 1718 2566 1721
rect 2670 1721 2673 1728
rect 2626 1718 2673 1721
rect 2690 1718 2702 1721
rect 2706 1718 3102 1721
rect 3170 1718 3310 1721
rect 3314 1718 3390 1721
rect 3434 1718 3438 1721
rect 3450 1718 3550 1721
rect 3738 1718 4110 1721
rect 4162 1718 4214 1721
rect 4222 1718 4230 1721
rect 4234 1718 4302 1721
rect 562 1708 702 1711
rect 922 1708 1102 1711
rect 1146 1708 1374 1711
rect 1394 1708 1574 1711
rect 1594 1708 1654 1711
rect 1918 1711 1921 1718
rect 1658 1708 1921 1711
rect 2010 1708 2022 1711
rect 2042 1708 2134 1711
rect 2138 1708 2273 1711
rect 2282 1708 2478 1711
rect 2482 1708 2574 1711
rect 2662 1708 2870 1711
rect 2874 1708 2918 1711
rect 2994 1708 2998 1711
rect 3034 1708 3054 1711
rect 3090 1708 3190 1711
rect 3202 1708 3286 1711
rect 3378 1708 3406 1711
rect 3418 1708 3542 1711
rect 3570 1708 3622 1711
rect 3650 1708 3678 1711
rect 3682 1708 3838 1711
rect 3890 1708 3902 1711
rect 3906 1708 3934 1711
rect 4002 1708 4062 1711
rect 4066 1708 4174 1711
rect 4234 1708 4246 1711
rect 896 1703 898 1707
rect 902 1703 905 1707
rect 910 1703 912 1707
rect 1928 1703 1930 1707
rect 1934 1703 1937 1707
rect 1942 1703 1944 1707
rect 818 1698 846 1701
rect 850 1698 889 1701
rect -26 1691 -22 1692
rect -26 1688 38 1691
rect 642 1688 678 1691
rect 746 1688 758 1691
rect 794 1688 798 1691
rect 886 1691 889 1698
rect 1426 1698 1494 1701
rect 1498 1698 1542 1701
rect 1546 1698 1598 1701
rect 1602 1698 1646 1701
rect 1658 1698 1830 1701
rect 1866 1698 1886 1701
rect 1962 1698 1998 1701
rect 2010 1698 2014 1701
rect 2050 1698 2054 1701
rect 2094 1698 2142 1701
rect 2178 1698 2238 1701
rect 2242 1698 2246 1701
rect 2270 1701 2273 1708
rect 2662 1701 2665 1708
rect 2952 1703 2954 1707
rect 2958 1703 2961 1707
rect 2966 1703 2968 1707
rect 2270 1698 2665 1701
rect 2706 1698 2710 1701
rect 2762 1698 2806 1701
rect 2842 1698 2862 1701
rect 2978 1698 3078 1701
rect 3082 1698 3174 1701
rect 3178 1698 3262 1701
rect 3266 1698 3302 1701
rect 3314 1698 3334 1701
rect 3418 1698 3510 1701
rect 3566 1701 3569 1708
rect 3976 1703 3978 1707
rect 3982 1703 3985 1707
rect 3990 1703 3992 1707
rect 3514 1698 3569 1701
rect 3706 1698 3718 1701
rect 3814 1698 3878 1701
rect 4106 1698 4318 1701
rect 886 1688 942 1691
rect 946 1688 966 1691
rect 974 1688 982 1691
rect 1138 1688 1302 1691
rect 1334 1691 1337 1698
rect 1334 1688 1342 1691
rect 1494 1688 1566 1691
rect 1570 1688 1622 1691
rect 1626 1688 1670 1691
rect 1754 1688 1790 1691
rect 1810 1688 1854 1691
rect 1910 1688 1918 1691
rect 1922 1688 1926 1691
rect 2094 1691 2097 1698
rect 1938 1688 2097 1691
rect 2102 1688 2110 1691
rect 2114 1688 2254 1691
rect 2266 1688 2278 1691
rect 2386 1688 2502 1691
rect 2590 1688 2686 1691
rect 2746 1688 2750 1691
rect 2770 1688 2774 1691
rect 2890 1688 3414 1691
rect 3450 1688 3454 1691
rect 3814 1691 3817 1698
rect 4358 1692 4361 1698
rect 3506 1688 3817 1691
rect 3826 1688 3830 1691
rect 4238 1688 4246 1691
rect 4250 1688 4350 1691
rect 170 1678 382 1681
rect 394 1678 502 1681
rect 770 1678 870 1681
rect 898 1678 1094 1681
rect 1106 1678 1174 1681
rect 1210 1678 1254 1681
rect 1282 1678 1286 1681
rect 1310 1681 1313 1688
rect 1306 1678 1313 1681
rect 1322 1678 1398 1681
rect 1414 1681 1417 1688
rect 1446 1682 1449 1688
rect 1494 1682 1497 1688
rect 1414 1678 1430 1681
rect 1554 1678 1574 1681
rect 1578 1678 1585 1681
rect 1634 1678 1654 1681
rect 1726 1681 1729 1688
rect 2590 1682 2593 1688
rect 1666 1678 1782 1681
rect 1786 1678 1822 1681
rect 1842 1678 1870 1681
rect 1874 1678 2014 1681
rect 2026 1678 2126 1681
rect 2402 1678 2590 1681
rect 2650 1678 2654 1681
rect 2782 1681 2785 1688
rect 2658 1678 2785 1681
rect 2830 1681 2833 1688
rect 2810 1678 2833 1681
rect 2930 1678 3166 1681
rect 3394 1678 3478 1681
rect 3498 1678 3510 1681
rect 3514 1678 3606 1681
rect 3610 1678 3622 1681
rect 3690 1678 3734 1681
rect 3754 1678 3758 1681
rect 3930 1678 4070 1681
rect 4082 1678 4222 1681
rect 4250 1678 4254 1681
rect 4274 1678 4374 1681
rect -26 1671 -22 1672
rect 6 1671 9 1678
rect -26 1668 9 1671
rect 158 1672 161 1678
rect 606 1672 609 1678
rect 718 1672 721 1678
rect 3070 1672 3073 1678
rect 346 1668 358 1671
rect 362 1668 422 1671
rect 478 1668 582 1671
rect 586 1668 590 1671
rect 730 1668 734 1671
rect 738 1668 758 1671
rect 762 1668 982 1671
rect 1018 1668 1038 1671
rect 1146 1668 1198 1671
rect 1250 1668 1366 1671
rect 1386 1668 1438 1671
rect 1442 1668 1454 1671
rect 1474 1668 1526 1671
rect 1538 1668 1686 1671
rect 1706 1668 1710 1671
rect 1722 1668 2121 1671
rect 2130 1668 2150 1671
rect 2154 1668 2161 1671
rect 2178 1668 2262 1671
rect 2586 1668 2846 1671
rect 3142 1668 3438 1671
rect 3442 1668 3518 1671
rect 3578 1668 3606 1671
rect 3610 1668 3617 1671
rect 3626 1668 4094 1671
rect 4114 1668 4166 1671
rect 4266 1668 4321 1671
rect 478 1662 481 1668
rect 34 1658 166 1661
rect 218 1658 246 1661
rect 386 1658 430 1661
rect 634 1658 814 1661
rect 818 1658 822 1661
rect 882 1658 902 1661
rect 914 1658 918 1661
rect 930 1658 934 1661
rect 962 1658 998 1661
rect 1050 1658 1214 1661
rect 1218 1658 1238 1661
rect 1242 1658 1374 1661
rect 1386 1658 1430 1661
rect 1458 1658 1462 1661
rect 1478 1658 1486 1661
rect 1490 1658 1502 1661
rect 1610 1658 1614 1661
rect 1698 1658 2022 1661
rect 2026 1658 2038 1661
rect 2066 1658 2086 1661
rect 2106 1658 2110 1661
rect 2118 1661 2121 1668
rect 2118 1658 2366 1661
rect 2370 1658 2398 1661
rect 2610 1658 2630 1661
rect 2658 1658 2718 1661
rect 3142 1661 3145 1668
rect 2762 1658 3145 1661
rect 3154 1658 3158 1661
rect 3162 1658 3206 1661
rect 3218 1658 3270 1661
rect 3274 1658 3406 1661
rect 3426 1658 3446 1661
rect 3530 1658 3614 1661
rect 3642 1658 3646 1661
rect 3682 1658 3734 1661
rect 3938 1658 3958 1661
rect 4010 1658 4030 1661
rect 4058 1658 4070 1661
rect 4114 1658 4134 1661
rect 4182 1661 4185 1668
rect 4198 1661 4201 1668
rect 4318 1662 4321 1668
rect 4182 1658 4201 1661
rect 4250 1658 4286 1661
rect 4342 1658 4358 1661
rect -26 1651 -22 1652
rect -26 1648 6 1651
rect 234 1648 254 1651
rect 258 1648 646 1651
rect 722 1648 742 1651
rect 754 1648 790 1651
rect 882 1648 950 1651
rect 1026 1648 1086 1651
rect 1090 1648 1102 1651
rect 1122 1648 1126 1651
rect 1218 1648 1233 1651
rect 1242 1648 1358 1651
rect 1370 1648 1390 1651
rect 1498 1648 1502 1651
rect 1510 1651 1513 1658
rect 1510 1648 1614 1651
rect 1650 1648 1750 1651
rect 1778 1648 1782 1651
rect 1786 1648 1790 1651
rect 1814 1648 1886 1651
rect 1914 1648 1918 1651
rect 1930 1648 1998 1651
rect 2010 1648 2070 1651
rect 2086 1651 2089 1658
rect 4342 1652 4345 1658
rect 2086 1648 2374 1651
rect 2506 1648 2606 1651
rect 2618 1648 2638 1651
rect 2714 1648 2718 1651
rect 2874 1648 3134 1651
rect 3186 1648 3190 1651
rect 3466 1648 3470 1651
rect 3518 1648 3550 1651
rect 3602 1648 3622 1651
rect 3690 1648 3694 1651
rect 3722 1648 3846 1651
rect 3946 1648 3950 1651
rect 4026 1648 4030 1651
rect 4050 1648 4078 1651
rect 4122 1648 4126 1651
rect 4146 1648 4150 1651
rect 4170 1648 4262 1651
rect 4290 1648 4294 1651
rect 4374 1651 4377 1658
rect 4370 1648 4377 1651
rect 974 1642 977 1648
rect 1230 1642 1233 1648
rect 1814 1642 1817 1648
rect 2830 1642 2833 1648
rect 3518 1642 3521 1648
rect 146 1638 310 1641
rect 314 1638 326 1641
rect 330 1638 398 1641
rect 506 1638 686 1641
rect 706 1638 710 1641
rect 714 1638 838 1641
rect 946 1638 958 1641
rect 978 1638 1038 1641
rect 1042 1638 1070 1641
rect 1098 1638 1190 1641
rect 1378 1638 1406 1641
rect 1466 1638 1590 1641
rect 1674 1638 1710 1641
rect 1714 1638 1758 1641
rect 1774 1638 1798 1641
rect 1866 1638 1942 1641
rect 1946 1638 2110 1641
rect 2138 1638 2142 1641
rect 2170 1638 2278 1641
rect 2594 1638 2662 1641
rect 2666 1638 2790 1641
rect 2850 1638 3182 1641
rect 3250 1638 3502 1641
rect 3662 1641 3665 1648
rect 3662 1638 3710 1641
rect 3946 1638 3966 1641
rect 4010 1638 4062 1641
rect 4122 1638 4142 1641
rect 4186 1638 4270 1641
rect 4338 1638 4366 1641
rect 686 1631 689 1638
rect 1262 1632 1265 1638
rect 1774 1632 1777 1638
rect 686 1628 838 1631
rect 874 1628 878 1631
rect 1010 1628 1150 1631
rect 1306 1628 1534 1631
rect 1538 1628 1582 1631
rect 1602 1628 1718 1631
rect 1866 1628 1961 1631
rect 1970 1628 1974 1631
rect 2002 1628 2198 1631
rect 2202 1628 2222 1631
rect 2626 1628 2742 1631
rect 2746 1628 3086 1631
rect 3130 1628 3254 1631
rect 3378 1628 3438 1631
rect 3442 1628 3606 1631
rect 3954 1628 4014 1631
rect 4018 1628 4046 1631
rect 4214 1628 4294 1631
rect 4314 1628 4342 1631
rect 1958 1622 1961 1628
rect 4214 1622 4217 1628
rect 4358 1622 4361 1628
rect 10 1618 417 1621
rect 666 1618 758 1621
rect 834 1618 1814 1621
rect 1842 1618 1854 1621
rect 1914 1618 1918 1621
rect 1970 1618 2062 1621
rect 2074 1618 2222 1621
rect 2602 1618 2646 1621
rect 2682 1618 2910 1621
rect 2970 1618 2974 1621
rect 2978 1618 2982 1621
rect 3130 1618 3998 1621
rect 4306 1618 4350 1621
rect 414 1611 417 1618
rect 414 1608 1062 1611
rect 1066 1608 1406 1611
rect 1578 1608 1622 1611
rect 1642 1608 1694 1611
rect 1698 1608 1774 1611
rect 1818 1608 1934 1611
rect 2090 1608 2094 1611
rect 2122 1608 2214 1611
rect 2570 1608 2678 1611
rect 3138 1608 3222 1611
rect 3274 1608 3382 1611
rect 3610 1608 3678 1611
rect 3842 1608 3886 1611
rect 4314 1608 4334 1611
rect 392 1603 394 1607
rect 398 1603 401 1607
rect 406 1603 408 1607
rect 1416 1603 1418 1607
rect 1422 1603 1425 1607
rect 1430 1603 1432 1607
rect 2440 1603 2442 1607
rect 2446 1603 2449 1607
rect 2454 1603 2456 1607
rect 3472 1603 3474 1607
rect 3478 1603 3481 1607
rect 3486 1603 3488 1607
rect 426 1598 638 1601
rect 642 1598 766 1601
rect 778 1598 886 1601
rect 1002 1598 1022 1601
rect 1106 1598 1166 1601
rect 1170 1598 1198 1601
rect 1238 1598 1278 1601
rect 1290 1598 1366 1601
rect 1370 1598 1390 1601
rect 1458 1598 1462 1601
rect 1474 1598 1542 1601
rect 1570 1598 1638 1601
rect 1658 1598 1990 1601
rect 2090 1598 2182 1601
rect 2290 1598 2422 1601
rect 2538 1598 2694 1601
rect 2722 1598 2878 1601
rect 2890 1598 3382 1601
rect 3642 1598 3678 1601
rect -26 1591 -22 1592
rect -26 1588 9 1591
rect 6 1582 9 1588
rect 322 1588 366 1591
rect 530 1588 697 1591
rect 714 1588 766 1591
rect 850 1588 854 1591
rect 902 1588 910 1591
rect 914 1588 1086 1591
rect 1122 1588 1134 1591
rect 1174 1588 1182 1591
rect 1238 1591 1241 1598
rect 1186 1588 1241 1591
rect 1410 1588 1518 1591
rect 1522 1588 1646 1591
rect 1666 1588 1950 1591
rect 1954 1588 2006 1591
rect 2014 1588 2022 1591
rect 2026 1588 2054 1591
rect 2058 1588 3126 1591
rect 3146 1588 3294 1591
rect 3418 1588 3494 1591
rect 3818 1588 3822 1591
rect 4038 1588 4222 1591
rect 4262 1588 4286 1591
rect 30 1581 33 1588
rect 694 1582 697 1588
rect 14 1578 33 1581
rect 330 1578 409 1581
rect 586 1578 606 1581
rect 718 1578 838 1581
rect 842 1578 878 1581
rect 890 1578 950 1581
rect 954 1578 958 1581
rect 1074 1578 1102 1581
rect 1110 1581 1113 1588
rect 1110 1578 1318 1581
rect 1322 1578 1326 1581
rect 1330 1578 1358 1581
rect 1498 1578 2734 1581
rect 2738 1578 2878 1581
rect 3186 1578 3262 1581
rect 3326 1581 3329 1588
rect 3290 1578 3329 1581
rect 3410 1578 3446 1581
rect 3466 1578 3582 1581
rect 3646 1581 3649 1588
rect 4038 1582 4041 1588
rect 4262 1582 4265 1588
rect 4326 1582 4329 1588
rect 3646 1578 3718 1581
rect 3722 1578 3790 1581
rect 3794 1578 3918 1581
rect 4274 1578 4326 1581
rect -26 1571 -22 1572
rect 14 1571 17 1578
rect -26 1568 17 1571
rect 126 1571 129 1578
rect 26 1568 129 1571
rect 146 1568 238 1571
rect 242 1568 398 1571
rect 406 1571 409 1578
rect 646 1571 649 1578
rect 406 1568 649 1571
rect 718 1571 721 1578
rect 698 1568 721 1571
rect 770 1568 774 1571
rect 778 1568 798 1571
rect 810 1568 814 1571
rect 842 1568 942 1571
rect 986 1568 1478 1571
rect 1530 1568 1566 1571
rect 1586 1568 1606 1571
rect 1618 1568 1630 1571
rect 1682 1568 1718 1571
rect 1778 1568 1838 1571
rect 1982 1568 2118 1571
rect 2274 1568 3166 1571
rect 3314 1568 3342 1571
rect 3402 1568 3470 1571
rect 3474 1568 3654 1571
rect 3658 1568 3662 1571
rect 3666 1568 3694 1571
rect 3698 1568 3702 1571
rect 4118 1571 4121 1578
rect 4118 1568 4142 1571
rect 4202 1568 4222 1571
rect 4322 1568 4326 1571
rect 90 1558 430 1561
rect 634 1558 678 1561
rect 726 1561 729 1568
rect 1982 1562 1985 1568
rect 2198 1562 2201 1568
rect 3294 1562 3297 1568
rect 3310 1562 3313 1568
rect 726 1558 742 1561
rect 746 1558 894 1561
rect 1034 1558 1070 1561
rect 1122 1558 1142 1561
rect 1146 1558 1190 1561
rect 1226 1558 1270 1561
rect 1282 1558 1302 1561
rect 1314 1558 1358 1561
rect 1434 1558 1502 1561
rect 1546 1558 1678 1561
rect 1726 1558 1734 1561
rect 1754 1558 1758 1561
rect 1762 1558 1790 1561
rect 1794 1558 1862 1561
rect 1954 1558 1969 1561
rect 2034 1558 2150 1561
rect 2154 1558 2158 1561
rect 2298 1558 2302 1561
rect 2362 1558 2550 1561
rect 2554 1558 2606 1561
rect 2614 1558 2638 1561
rect 2690 1558 2726 1561
rect 2738 1558 2822 1561
rect 2842 1558 2886 1561
rect 2890 1558 3142 1561
rect 3250 1558 3270 1561
rect 3330 1558 3334 1561
rect 3338 1558 3366 1561
rect 3466 1558 3622 1561
rect 3630 1558 3638 1561
rect 3642 1558 3670 1561
rect 3690 1558 3782 1561
rect 3862 1561 3865 1568
rect 3842 1558 3865 1561
rect 3886 1562 3889 1568
rect 3930 1558 3934 1561
rect 3946 1558 3990 1561
rect 4042 1558 4046 1561
rect 4090 1558 4102 1561
rect 4146 1558 4190 1561
rect 4194 1558 4246 1561
rect 1510 1552 1513 1558
rect -26 1551 -22 1552
rect -26 1548 14 1551
rect 74 1548 134 1551
rect 138 1548 174 1551
rect 178 1548 430 1551
rect 770 1548 814 1551
rect 866 1548 870 1551
rect 898 1548 902 1551
rect 970 1548 974 1551
rect 1010 1548 1022 1551
rect 1058 1548 1086 1551
rect 1098 1548 1150 1551
rect 1258 1548 1462 1551
rect 1554 1548 1558 1551
rect 1678 1551 1681 1558
rect 1666 1548 1681 1551
rect 1726 1552 1729 1558
rect 1966 1552 1969 1558
rect 1998 1552 2001 1558
rect 2614 1552 2617 1558
rect 1810 1548 1814 1551
rect 1842 1548 1870 1551
rect 1898 1548 1902 1551
rect 2122 1548 2158 1551
rect 2186 1548 2246 1551
rect 2442 1548 2558 1551
rect 2562 1548 2569 1551
rect 2578 1548 2582 1551
rect 2626 1548 2654 1551
rect 2674 1548 2710 1551
rect 2722 1548 2782 1551
rect 2786 1548 2822 1551
rect 2890 1548 2894 1551
rect 2946 1548 2982 1551
rect 3138 1548 3166 1551
rect 3174 1551 3177 1558
rect 3206 1551 3209 1558
rect 3398 1552 3401 1558
rect 3414 1552 3417 1558
rect 3174 1548 3209 1551
rect 3218 1548 3326 1551
rect 3330 1548 3374 1551
rect 3434 1548 3462 1551
rect 3554 1548 3558 1551
rect 3578 1548 3638 1551
rect 3822 1551 3825 1558
rect 3642 1548 3825 1551
rect 3842 1548 3902 1551
rect 3906 1548 4206 1551
rect 4250 1548 4270 1551
rect 4298 1548 4310 1551
rect 1654 1542 1657 1548
rect 1798 1542 1801 1548
rect 1830 1542 1833 1548
rect 106 1538 142 1541
rect 226 1538 310 1541
rect 386 1538 478 1541
rect 618 1538 670 1541
rect 690 1538 694 1541
rect 698 1538 718 1541
rect 842 1538 926 1541
rect 966 1538 1014 1541
rect 1058 1538 1126 1541
rect 1298 1538 1438 1541
rect 1482 1538 1486 1541
rect 1490 1538 1550 1541
rect 1618 1538 1630 1541
rect 1682 1538 1750 1541
rect 1842 1538 1894 1541
rect 1946 1538 1958 1541
rect 2026 1538 2094 1541
rect 2106 1538 2118 1541
rect 2266 1538 2366 1541
rect 2370 1538 2374 1541
rect 2474 1538 2750 1541
rect 2754 1538 3070 1541
rect 3574 1541 3577 1548
rect 3074 1538 3577 1541
rect 3586 1538 3590 1541
rect 3626 1538 3630 1541
rect 3722 1538 3734 1541
rect 3762 1538 3766 1541
rect 3802 1538 3918 1541
rect 3930 1538 3934 1541
rect 4002 1538 4102 1541
rect 4170 1538 4174 1541
rect 4186 1538 4214 1541
rect 4230 1541 4233 1548
rect 4230 1538 4246 1541
rect 870 1532 873 1538
rect 966 1532 969 1538
rect 1262 1532 1265 1538
rect 1446 1532 1449 1538
rect -26 1531 -22 1532
rect -26 1528 198 1531
rect 578 1528 638 1531
rect 642 1528 742 1531
rect 1138 1528 1214 1531
rect 1218 1528 1257 1531
rect 1274 1528 1334 1531
rect 1362 1528 1369 1531
rect 1450 1528 1582 1531
rect 1586 1528 1590 1531
rect 1926 1531 1929 1538
rect 2422 1532 2425 1538
rect 3686 1532 3689 1538
rect 1634 1528 1929 1531
rect 1994 1528 2134 1531
rect 2138 1528 2174 1531
rect 2178 1528 2182 1531
rect 2210 1528 2422 1531
rect 2490 1528 2526 1531
rect 2594 1528 2598 1531
rect 2642 1528 2670 1531
rect 2786 1528 2790 1531
rect 3146 1528 3150 1531
rect 3158 1528 3166 1531
rect 3186 1528 3190 1531
rect 3202 1528 3206 1531
rect 3254 1528 3278 1531
rect 3302 1528 3318 1531
rect 3338 1528 3342 1531
rect 3362 1528 3366 1531
rect 3378 1528 3454 1531
rect 3458 1528 3502 1531
rect 3514 1528 3518 1531
rect 3530 1528 3534 1531
rect 3546 1528 3574 1531
rect 3586 1528 3590 1531
rect 3626 1528 3654 1531
rect 3706 1528 3742 1531
rect 3778 1528 3958 1531
rect 4162 1528 4342 1531
rect 170 1518 422 1521
rect 490 1518 838 1521
rect 874 1518 1006 1521
rect 1010 1518 1046 1521
rect 1082 1518 1134 1521
rect 1138 1518 1238 1521
rect 1254 1521 1257 1528
rect 1366 1522 1369 1528
rect 3054 1522 3057 1528
rect 3158 1522 3161 1528
rect 3254 1522 3257 1528
rect 3302 1522 3305 1528
rect 3350 1522 3353 1528
rect 3374 1522 3377 1528
rect 1254 1518 1286 1521
rect 1442 1518 1606 1521
rect 1898 1518 1958 1521
rect 1978 1518 2046 1521
rect 2138 1518 2262 1521
rect 2346 1518 2350 1521
rect 2426 1518 2510 1521
rect 2562 1518 2598 1521
rect 2602 1518 2630 1521
rect 2746 1518 2846 1521
rect 2946 1518 2982 1521
rect 2986 1518 3054 1521
rect 3170 1518 3254 1521
rect 3418 1518 3430 1521
rect 3442 1518 3470 1521
rect 3498 1518 3502 1521
rect 3538 1518 3558 1521
rect 3598 1521 3601 1528
rect 3598 1518 3718 1521
rect 3730 1518 3814 1521
rect 3818 1518 3854 1521
rect 3946 1518 4054 1521
rect 4170 1518 4286 1521
rect -26 1508 -22 1512
rect 10 1508 870 1511
rect 962 1508 990 1511
rect 1202 1508 1294 1511
rect 1346 1508 1366 1511
rect 1394 1508 1406 1511
rect 1450 1508 1622 1511
rect 1642 1508 1686 1511
rect 1714 1508 1726 1511
rect 1794 1508 1846 1511
rect 1850 1508 1910 1511
rect 1978 1508 2070 1511
rect 2306 1508 2718 1511
rect 2874 1508 2910 1511
rect 2914 1508 2926 1511
rect 3042 1508 3462 1511
rect 3482 1508 3574 1511
rect 3618 1508 3654 1511
rect 3722 1508 3742 1511
rect 3746 1508 3750 1511
rect 3850 1508 3902 1511
rect 4050 1508 4062 1511
rect -26 1501 -23 1508
rect 896 1503 898 1507
rect 902 1503 905 1507
rect 910 1503 912 1507
rect 1928 1503 1930 1507
rect 1934 1503 1937 1507
rect 1942 1503 1944 1507
rect 2952 1503 2954 1507
rect 2958 1503 2961 1507
rect 2966 1503 2968 1507
rect 3976 1503 3978 1507
rect 3982 1503 3985 1507
rect 3990 1503 3992 1507
rect -26 1498 6 1501
rect 42 1498 78 1501
rect 82 1498 358 1501
rect 618 1498 782 1501
rect 786 1498 814 1501
rect 842 1498 846 1501
rect 858 1498 886 1501
rect 986 1498 1014 1501
rect 1210 1498 1342 1501
rect 1354 1498 1409 1501
rect 1466 1498 1470 1501
rect 1626 1498 1670 1501
rect 1690 1498 1734 1501
rect 2042 1498 2246 1501
rect 2338 1498 2558 1501
rect 2562 1498 2654 1501
rect 2658 1498 2686 1501
rect 2978 1498 3222 1501
rect 3242 1498 3302 1501
rect 3394 1498 3422 1501
rect 3438 1498 3969 1501
rect 4010 1498 4014 1501
rect 4018 1498 4070 1501
rect 4074 1498 4238 1501
rect -26 1491 -22 1492
rect -26 1488 6 1491
rect 18 1488 926 1491
rect 930 1488 1046 1491
rect 1050 1488 1062 1491
rect 1066 1488 1070 1491
rect 1074 1488 1182 1491
rect 1194 1488 1222 1491
rect 1330 1488 1390 1491
rect 1406 1491 1409 1498
rect 3438 1492 3441 1498
rect 1406 1488 1470 1491
rect 1474 1488 1481 1491
rect 1490 1488 1678 1491
rect 1714 1488 1766 1491
rect 1786 1488 1974 1491
rect 2234 1488 2382 1491
rect 2410 1488 2558 1491
rect 2570 1488 2606 1491
rect 2714 1488 2774 1491
rect 2802 1488 2814 1491
rect 2818 1488 2982 1491
rect 3102 1488 3318 1491
rect 3322 1488 3438 1491
rect 3554 1488 3606 1491
rect 3610 1488 3630 1491
rect 3770 1488 3798 1491
rect 3966 1491 3969 1498
rect 3966 1488 4206 1491
rect 34 1478 62 1481
rect 66 1478 78 1481
rect 274 1478 302 1481
rect 486 1478 518 1481
rect 570 1478 670 1481
rect 722 1478 801 1481
rect 834 1478 838 1481
rect 842 1478 1310 1481
rect 1398 1481 1401 1488
rect 1362 1478 1401 1481
rect 1418 1478 1518 1481
rect 1530 1478 1534 1481
rect 1686 1481 1689 1488
rect 3102 1482 3105 1488
rect 1674 1478 1689 1481
rect 1706 1478 1710 1481
rect 1754 1478 1758 1481
rect 1826 1478 1838 1481
rect 1890 1478 1926 1481
rect 2194 1478 2217 1481
rect -26 1471 -22 1472
rect -26 1468 6 1471
rect 50 1468 54 1471
rect 82 1468 166 1471
rect 182 1461 185 1478
rect 350 1471 353 1478
rect 486 1472 489 1478
rect 798 1472 801 1478
rect 2214 1472 2217 1478
rect 2514 1478 2694 1481
rect 2706 1478 2734 1481
rect 2834 1478 2838 1481
rect 3282 1478 3302 1481
rect 3322 1478 3334 1481
rect 3354 1478 3358 1481
rect 3386 1478 3422 1481
rect 3534 1481 3537 1488
rect 3710 1482 3713 1488
rect 3734 1482 3737 1488
rect 3942 1482 3945 1488
rect 3534 1478 3558 1481
rect 3562 1478 3606 1481
rect 3682 1478 3710 1481
rect 3738 1478 3782 1481
rect 3794 1478 3830 1481
rect 4066 1478 4129 1481
rect 4138 1478 4158 1481
rect 4162 1478 4198 1481
rect 4310 1481 4313 1488
rect 4218 1478 4313 1481
rect 350 1468 414 1471
rect 538 1468 630 1471
rect 650 1468 654 1471
rect 658 1468 726 1471
rect 754 1468 758 1471
rect 818 1468 878 1471
rect 890 1468 902 1471
rect 906 1468 974 1471
rect 978 1468 1086 1471
rect 1370 1468 1446 1471
rect 1498 1468 1502 1471
rect 1530 1468 1574 1471
rect 1762 1468 1774 1471
rect 1818 1468 1830 1471
rect 1898 1468 1902 1471
rect 2074 1468 2118 1471
rect 2230 1471 2233 1478
rect 3222 1472 3225 1478
rect 2230 1468 2326 1471
rect 2410 1468 2454 1471
rect 2458 1468 2478 1471
rect 2582 1468 2678 1471
rect 2730 1468 2750 1471
rect 2786 1468 2806 1471
rect 2810 1468 2830 1471
rect 3034 1468 3086 1471
rect 3106 1468 3110 1471
rect 3298 1468 3302 1471
rect 3330 1468 3334 1471
rect 3346 1468 3358 1471
rect 3370 1468 3374 1471
rect 3410 1468 3414 1471
rect 3434 1468 3470 1471
rect 3514 1468 3566 1471
rect 3570 1468 3590 1471
rect 3594 1468 3622 1471
rect 3642 1468 3694 1471
rect 3802 1468 3806 1471
rect 4126 1471 4129 1478
rect 4126 1468 4142 1471
rect 4194 1468 4238 1471
rect 4274 1468 4278 1471
rect 4306 1468 4310 1471
rect 510 1462 513 1468
rect 182 1458 502 1461
rect 602 1458 606 1461
rect 626 1458 638 1461
rect 658 1458 726 1461
rect 754 1458 774 1461
rect 794 1458 958 1461
rect 994 1458 1006 1461
rect 1126 1458 1142 1461
rect 1258 1458 1289 1461
rect 1346 1458 1358 1461
rect 1410 1458 1510 1461
rect 1570 1458 1574 1461
rect 1586 1458 1590 1461
rect 1598 1461 1601 1468
rect 1686 1462 1689 1468
rect 2390 1462 2393 1468
rect 2582 1462 2585 1468
rect 1598 1458 1654 1461
rect 1754 1458 1782 1461
rect 1786 1458 1822 1461
rect 1858 1458 1910 1461
rect 1946 1458 1974 1461
rect 2002 1458 2014 1461
rect 2114 1458 2302 1461
rect 2310 1458 2334 1461
rect 2338 1458 2374 1461
rect 2394 1458 2422 1461
rect 2642 1458 2718 1461
rect 2730 1458 2793 1461
rect 2826 1458 2830 1461
rect 2846 1461 2849 1468
rect 2846 1458 2870 1461
rect 2874 1458 2878 1461
rect 2898 1458 2902 1461
rect 3058 1458 3126 1461
rect 3130 1458 3166 1461
rect 3282 1458 3574 1461
rect 3578 1458 3838 1461
rect 3842 1458 3894 1461
rect 4058 1458 4086 1461
rect 4102 1461 4105 1468
rect 4118 1461 4121 1468
rect 4102 1458 4121 1461
rect 4170 1458 4230 1461
rect 4242 1458 4302 1461
rect 4306 1458 4318 1461
rect -26 1451 -22 1452
rect -26 1448 78 1451
rect 506 1448 566 1451
rect 610 1448 878 1451
rect 882 1448 982 1451
rect 986 1448 1038 1451
rect 1054 1451 1057 1458
rect 1042 1448 1057 1451
rect 1126 1452 1129 1458
rect 1286 1452 1289 1458
rect 2310 1452 2313 1458
rect 2790 1452 2793 1458
rect 4086 1452 4089 1458
rect 1322 1448 1390 1451
rect 1450 1448 1454 1451
rect 1458 1448 1470 1451
rect 1650 1448 1654 1451
rect 1666 1448 1782 1451
rect 1794 1448 1798 1451
rect 1834 1448 1870 1451
rect 1874 1448 2006 1451
rect 2054 1448 2062 1451
rect 2066 1448 2094 1451
rect 2362 1448 2398 1451
rect 2418 1448 2422 1451
rect 2482 1448 2654 1451
rect 2658 1448 2734 1451
rect 2754 1448 2766 1451
rect 3086 1448 3094 1451
rect 3098 1448 3318 1451
rect 3338 1448 3350 1451
rect 3362 1448 3393 1451
rect 3418 1448 3446 1451
rect 3554 1448 3670 1451
rect 3682 1448 3822 1451
rect 3826 1448 3854 1451
rect 3954 1448 4081 1451
rect 4114 1448 4166 1451
rect 4290 1448 4374 1451
rect 458 1438 518 1441
rect 554 1438 558 1441
rect 562 1438 590 1441
rect 682 1438 694 1441
rect 698 1438 790 1441
rect 802 1438 918 1441
rect 922 1438 966 1441
rect 1006 1438 1014 1441
rect 1018 1438 1022 1441
rect 1026 1438 1118 1441
rect 1386 1438 1406 1441
rect 1426 1438 1438 1441
rect 1442 1438 1502 1441
rect 1510 1441 1513 1448
rect 1510 1438 1670 1441
rect 1706 1438 1870 1441
rect 1914 1438 1990 1441
rect 2022 1441 2025 1448
rect 3390 1442 3393 1448
rect 4078 1442 4081 1448
rect 2022 1438 2214 1441
rect 2498 1438 3382 1441
rect 3410 1438 3414 1441
rect 3634 1438 3646 1441
rect 3650 1438 3678 1441
rect 3762 1438 3790 1441
rect 3794 1438 3910 1441
rect 3946 1438 4062 1441
rect 4106 1438 4150 1441
rect 4202 1438 4214 1441
rect 534 1431 537 1438
rect 442 1428 537 1431
rect 554 1428 598 1431
rect 650 1428 686 1431
rect 714 1428 822 1431
rect 826 1428 846 1431
rect 874 1428 1270 1431
rect 1282 1428 1686 1431
rect 1690 1428 2126 1431
rect 2314 1428 2438 1431
rect 2442 1428 2814 1431
rect 2890 1428 3430 1431
rect 3434 1428 3550 1431
rect 3586 1428 3598 1431
rect 3602 1428 3734 1431
rect 4090 1428 4182 1431
rect 4342 1431 4345 1438
rect 4226 1428 4345 1431
rect 10 1418 686 1421
rect 698 1418 806 1421
rect 890 1418 1078 1421
rect 1082 1418 1158 1421
rect 1162 1418 1974 1421
rect 2098 1418 2382 1421
rect 2430 1418 2438 1421
rect 2442 1418 2510 1421
rect 2530 1418 2710 1421
rect 2714 1418 2734 1421
rect 2838 1421 2841 1428
rect 2738 1418 2841 1421
rect 2858 1418 3374 1421
rect 3378 1418 3438 1421
rect 3442 1418 3454 1421
rect 3586 1418 3598 1421
rect 3626 1418 3854 1421
rect 4194 1418 4262 1421
rect 4330 1418 4350 1421
rect 418 1408 758 1411
rect 786 1408 862 1411
rect 898 1408 1006 1411
rect 1186 1408 1302 1411
rect 1378 1408 1406 1411
rect 1442 1408 1558 1411
rect 1578 1408 2262 1411
rect 2594 1408 2670 1411
rect 2674 1408 2718 1411
rect 2722 1408 2742 1411
rect 2746 1408 2886 1411
rect 2890 1408 3086 1411
rect 3090 1408 3462 1411
rect 3730 1408 3742 1411
rect 3914 1408 4022 1411
rect 392 1403 394 1407
rect 398 1403 401 1407
rect 406 1403 408 1407
rect 1416 1403 1418 1407
rect 1422 1403 1425 1407
rect 1430 1403 1432 1407
rect 2440 1403 2442 1407
rect 2446 1403 2449 1407
rect 2454 1403 2456 1407
rect 138 1398 342 1401
rect 538 1398 574 1401
rect 578 1398 606 1401
rect 610 1398 766 1401
rect 770 1398 806 1401
rect 810 1398 870 1401
rect 1194 1398 1206 1401
rect 1218 1398 1318 1401
rect 1474 1398 1590 1401
rect 1594 1398 1638 1401
rect 1642 1398 1654 1401
rect 1658 1398 1854 1401
rect 1922 1398 2038 1401
rect 2466 1398 2526 1401
rect 2590 1401 2593 1408
rect 3472 1403 3474 1407
rect 3478 1403 3481 1407
rect 3486 1403 3488 1407
rect 2570 1398 2593 1401
rect 2850 1398 2934 1401
rect 2938 1398 2974 1401
rect 3002 1398 3046 1401
rect 3098 1398 3366 1401
rect 3498 1398 3806 1401
rect 3906 1398 3934 1401
rect 3938 1398 4222 1401
rect -26 1391 -22 1392
rect -26 1388 94 1391
rect 186 1388 254 1391
rect 362 1388 486 1391
rect 690 1388 1182 1391
rect 1274 1388 1342 1391
rect 1394 1388 1505 1391
rect 1610 1388 1670 1391
rect 1722 1388 1726 1391
rect 1754 1388 1774 1391
rect 1850 1388 1878 1391
rect 1902 1388 1918 1391
rect 2010 1388 2038 1391
rect 2346 1388 2350 1391
rect 2386 1388 2438 1391
rect 2474 1388 2494 1391
rect 2514 1388 2550 1391
rect 2618 1388 2838 1391
rect 2850 1388 3278 1391
rect 3394 1388 3526 1391
rect 4182 1388 4190 1391
rect 4194 1388 4230 1391
rect 1502 1382 1505 1388
rect 1902 1382 1905 1388
rect 106 1378 142 1381
rect 354 1378 470 1381
rect 754 1378 798 1381
rect 850 1378 1190 1381
rect 1202 1378 1390 1381
rect 1418 1378 1462 1381
rect 1482 1378 1494 1381
rect 1562 1378 1638 1381
rect 1650 1378 1718 1381
rect 1722 1378 1726 1381
rect 1982 1381 1985 1388
rect 1982 1378 2046 1381
rect 2050 1378 2102 1381
rect 2114 1378 2118 1381
rect 2290 1378 2318 1381
rect 2358 1381 2361 1388
rect 2358 1378 2478 1381
rect 2482 1378 2486 1381
rect 2494 1378 2502 1381
rect 2506 1378 2558 1381
rect 2562 1378 2630 1381
rect 2634 1378 2726 1381
rect 2730 1378 3950 1381
rect 3962 1378 4038 1381
rect 4042 1378 4070 1381
rect 4074 1378 4086 1381
rect 4090 1378 4134 1381
rect 4138 1378 4166 1381
rect 4170 1378 4374 1381
rect -26 1371 -22 1372
rect 6 1371 9 1378
rect -26 1368 9 1371
rect 62 1371 65 1378
rect 50 1368 65 1371
rect 82 1368 670 1371
rect 802 1368 854 1371
rect 1010 1368 1046 1371
rect 1226 1368 1958 1371
rect 1962 1368 2630 1371
rect 2794 1368 2814 1371
rect 2834 1368 3030 1371
rect 3202 1368 3318 1371
rect 3386 1368 3526 1371
rect 3546 1368 3697 1371
rect 3706 1368 3838 1371
rect 3978 1368 4038 1371
rect 4042 1368 4049 1371
rect 4058 1368 4062 1371
rect 4082 1368 4150 1371
rect 4154 1368 4182 1371
rect 4218 1368 4286 1371
rect 26 1358 126 1361
rect 234 1358 366 1361
rect 562 1358 729 1361
rect 738 1358 846 1361
rect 866 1358 902 1361
rect 914 1358 918 1361
rect 942 1361 945 1368
rect 3694 1362 3697 1368
rect 4046 1362 4049 1368
rect 930 1358 945 1361
rect 1050 1358 1078 1361
rect 1162 1358 1246 1361
rect 1298 1358 1326 1361
rect 1338 1358 1342 1361
rect 1354 1358 1358 1361
rect 1378 1358 1422 1361
rect 1450 1358 1550 1361
rect 1626 1358 1630 1361
rect 1650 1358 1758 1361
rect 1770 1358 1838 1361
rect 1878 1358 1886 1361
rect 1962 1358 1966 1361
rect 2010 1358 2014 1361
rect 2026 1358 2054 1361
rect 2066 1358 2070 1361
rect 2106 1358 2302 1361
rect 2322 1358 2326 1361
rect 2402 1358 2422 1361
rect 2430 1358 2526 1361
rect 2586 1358 2590 1361
rect 2666 1358 2686 1361
rect 2794 1358 2806 1361
rect 2810 1358 3070 1361
rect 3218 1358 3230 1361
rect 3334 1358 3342 1361
rect 3346 1358 3542 1361
rect 3746 1358 3750 1361
rect 3778 1358 3782 1361
rect 4018 1358 4022 1361
rect 4050 1358 4094 1361
rect 4122 1358 4126 1361
rect 4290 1358 4294 1361
rect 4298 1358 4334 1361
rect -26 1351 -22 1352
rect -26 1348 30 1351
rect 58 1348 110 1351
rect 114 1348 126 1351
rect 306 1348 374 1351
rect 498 1348 518 1351
rect 706 1348 710 1351
rect 726 1351 729 1358
rect 726 1348 790 1351
rect 810 1348 830 1351
rect 842 1348 918 1351
rect 1058 1348 1062 1351
rect 1074 1348 1094 1351
rect 1150 1351 1153 1358
rect 1150 1348 1174 1351
rect 1194 1348 1230 1351
rect 1266 1348 1270 1351
rect 1306 1348 1318 1351
rect 1322 1348 1446 1351
rect 1450 1348 1454 1351
rect 1482 1348 1486 1351
rect 1530 1348 1630 1351
rect 1682 1348 1694 1351
rect 1738 1348 1742 1351
rect 1762 1348 1766 1351
rect 1778 1348 1814 1351
rect 1818 1348 1846 1351
rect 1858 1348 1870 1351
rect 1890 1348 1894 1351
rect 1962 1348 2286 1351
rect 2318 1351 2321 1358
rect 2306 1348 2321 1351
rect 2338 1348 2342 1351
rect 2354 1348 2390 1351
rect 2430 1351 2433 1358
rect 2410 1348 2433 1351
rect 2490 1348 2494 1351
rect 2574 1351 2577 1358
rect 2554 1348 2577 1351
rect 2622 1351 2625 1358
rect 3270 1352 3273 1358
rect 2622 1348 2654 1351
rect 2690 1348 2718 1351
rect 2778 1348 2806 1351
rect 2930 1348 2950 1351
rect 3018 1348 3022 1351
rect 3234 1348 3262 1351
rect 3282 1348 3398 1351
rect 3610 1348 3614 1351
rect 3618 1348 3710 1351
rect 3714 1348 3790 1351
rect 3806 1351 3809 1358
rect 3830 1351 3833 1358
rect 4150 1352 4153 1358
rect 3806 1348 3870 1351
rect 3938 1348 3950 1351
rect 3970 1348 3990 1351
rect 4026 1348 4094 1351
rect 4122 1348 4126 1351
rect 4186 1348 4254 1351
rect 4258 1348 4342 1351
rect 58 1338 102 1341
rect 682 1338 710 1341
rect 722 1338 750 1341
rect 866 1338 886 1341
rect 898 1338 942 1341
rect 946 1338 1014 1341
rect 1042 1338 1118 1341
rect 1122 1338 1134 1341
rect 1154 1338 1166 1341
rect 1226 1338 1230 1341
rect 1298 1338 1302 1341
rect 1370 1338 1374 1341
rect 1402 1338 1478 1341
rect 1554 1338 1574 1341
rect 1586 1338 1902 1341
rect 1914 1338 1990 1341
rect 2298 1338 2742 1341
rect 2746 1338 2798 1341
rect 2818 1338 2862 1341
rect 2866 1338 2934 1341
rect 2938 1338 3014 1341
rect 3166 1338 3174 1341
rect 3250 1338 3254 1341
rect 3306 1338 3310 1341
rect 3346 1338 3350 1341
rect 3370 1338 3598 1341
rect 3610 1338 3638 1341
rect 3650 1338 3654 1341
rect 3666 1338 3670 1341
rect 3674 1338 3878 1341
rect 3882 1338 4206 1341
rect 4218 1338 4302 1341
rect 4314 1338 4358 1341
rect 246 1332 249 1338
rect 2054 1332 2057 1338
rect 3166 1332 3169 1338
rect 3286 1332 3289 1338
rect 578 1328 742 1331
rect 762 1328 838 1331
rect 846 1328 1054 1331
rect 1146 1328 1414 1331
rect 1426 1328 1838 1331
rect 1842 1328 1926 1331
rect 1954 1328 1998 1331
rect 2378 1328 2398 1331
rect 2434 1328 2526 1331
rect 2530 1328 2598 1331
rect 2602 1328 2606 1331
rect 2642 1328 2654 1331
rect 2714 1328 2750 1331
rect 2842 1328 2846 1331
rect 2858 1328 2894 1331
rect 2970 1328 3038 1331
rect 3294 1331 3297 1338
rect 3294 1328 3318 1331
rect 3330 1328 3334 1331
rect 3346 1328 3358 1331
rect 3362 1328 3438 1331
rect 3530 1328 3542 1331
rect 3562 1328 3654 1331
rect 3674 1328 3694 1331
rect 3786 1328 3918 1331
rect 4010 1328 4030 1331
rect 4034 1328 4110 1331
rect 4114 1328 4126 1331
rect 4178 1328 4190 1331
rect 4258 1328 4318 1331
rect 482 1318 662 1321
rect 666 1318 742 1321
rect 846 1321 849 1328
rect 2622 1322 2625 1328
rect 762 1318 849 1321
rect 930 1318 934 1321
rect 938 1318 1054 1321
rect 1078 1318 1230 1321
rect 1250 1318 1294 1321
rect 1330 1318 1462 1321
rect 1478 1318 1486 1321
rect 1610 1318 1614 1321
rect 1634 1318 1638 1321
rect 1698 1318 1702 1321
rect 1730 1318 1734 1321
rect 1746 1318 1750 1321
rect 1770 1318 1782 1321
rect 1802 1318 1806 1321
rect 1858 1318 1870 1321
rect 1882 1318 1886 1321
rect 1894 1318 2102 1321
rect 2154 1318 2158 1321
rect 2202 1318 2406 1321
rect 2630 1318 3734 1321
rect 3738 1318 3798 1321
rect 4234 1318 4254 1321
rect 4266 1318 4286 1321
rect 466 1308 694 1311
rect 754 1308 766 1311
rect 770 1308 822 1311
rect 970 1308 974 1311
rect 1078 1311 1081 1318
rect 1566 1312 1569 1318
rect 1574 1312 1577 1318
rect 1026 1308 1081 1311
rect 1090 1308 1390 1311
rect 1474 1308 1486 1311
rect 1514 1308 1542 1311
rect 1594 1308 1710 1311
rect 1738 1308 1830 1311
rect 1894 1311 1897 1318
rect 1890 1308 1897 1311
rect 2034 1308 2078 1311
rect 2082 1308 2086 1311
rect 2630 1311 2633 1318
rect 2098 1308 2633 1311
rect 2642 1308 2670 1311
rect 2674 1308 2870 1311
rect 3026 1308 3902 1311
rect 4186 1308 4238 1311
rect 4250 1308 4262 1311
rect 4386 1308 4390 1311
rect 896 1303 898 1307
rect 902 1303 905 1307
rect 910 1303 912 1307
rect 1928 1303 1930 1307
rect 1934 1303 1937 1307
rect 1942 1303 1944 1307
rect 2952 1303 2954 1307
rect 2958 1303 2961 1307
rect 2966 1303 2968 1307
rect 3976 1303 3978 1307
rect 3982 1303 3985 1307
rect 3990 1303 3992 1307
rect -26 1301 -22 1302
rect -26 1298 6 1301
rect 218 1298 422 1301
rect 690 1298 718 1301
rect 794 1298 854 1301
rect 962 1298 974 1301
rect 1018 1298 1166 1301
rect 1170 1298 1382 1301
rect 1394 1298 1526 1301
rect 1538 1298 1686 1301
rect 1690 1298 1790 1301
rect 1794 1298 1814 1301
rect 1818 1298 1894 1301
rect 2074 1298 2526 1301
rect 2538 1298 2753 1301
rect 3034 1298 3150 1301
rect 3266 1298 3294 1301
rect 3382 1298 3414 1301
rect 3434 1298 3454 1301
rect 3482 1298 3806 1301
rect 4106 1298 4118 1301
rect 4246 1301 4249 1308
rect 4122 1298 4249 1301
rect 266 1288 590 1291
rect 666 1288 774 1291
rect 826 1288 886 1291
rect 946 1288 1070 1291
rect 1082 1288 1094 1291
rect 1114 1288 1198 1291
rect 1346 1288 1350 1291
rect 1358 1288 1366 1291
rect 1370 1288 1814 1291
rect 1818 1288 2038 1291
rect 2634 1288 2726 1291
rect 2750 1291 2753 1298
rect 2750 1288 2974 1291
rect 3066 1288 3070 1291
rect 3074 1288 3134 1291
rect 3142 1288 3150 1291
rect 3154 1288 3174 1291
rect 3178 1288 3222 1291
rect 3382 1291 3385 1298
rect 3242 1288 3385 1291
rect 3426 1288 3430 1291
rect 3506 1288 3534 1291
rect 3538 1288 3614 1291
rect 3706 1288 3726 1291
rect 3730 1288 3742 1291
rect 3754 1288 3758 1291
rect 3762 1288 3798 1291
rect 3818 1288 3862 1291
rect 3898 1288 3910 1291
rect 3914 1288 3926 1291
rect 3930 1288 3942 1291
rect 3946 1288 4214 1291
rect -26 1281 -22 1282
rect -26 1278 14 1281
rect 94 1278 142 1281
rect 262 1281 265 1288
rect 146 1278 265 1281
rect 518 1278 550 1281
rect 554 1278 558 1281
rect 594 1278 702 1281
rect 730 1278 998 1281
rect 1090 1278 1102 1281
rect 1130 1278 1134 1281
rect 1186 1278 1206 1281
rect 1230 1281 1233 1288
rect 2062 1282 2065 1288
rect 1230 1278 1286 1281
rect 1290 1278 1366 1281
rect 1370 1278 1398 1281
rect 1402 1278 1534 1281
rect 1546 1278 1769 1281
rect 94 1272 97 1278
rect 518 1272 521 1278
rect 1766 1272 1769 1278
rect 1882 1278 1990 1281
rect 1994 1278 2014 1281
rect 2226 1278 2286 1281
rect 2290 1278 2294 1281
rect 2518 1281 2521 1288
rect 2742 1282 2745 1288
rect 3686 1282 3689 1288
rect 3878 1282 3881 1288
rect 2518 1278 2694 1281
rect 2698 1278 2734 1281
rect 2802 1278 2806 1281
rect 2810 1278 2822 1281
rect 2994 1278 3046 1281
rect 3050 1278 3126 1281
rect 3130 1278 3166 1281
rect 3178 1278 3310 1281
rect 3330 1278 3358 1281
rect 3362 1278 3382 1281
rect 3394 1278 3398 1281
rect 3422 1278 3462 1281
rect 3658 1278 3678 1281
rect 3698 1278 3782 1281
rect 3786 1278 3822 1281
rect 3922 1278 4086 1281
rect 4122 1278 4198 1281
rect 4202 1278 4286 1281
rect 4338 1278 4374 1281
rect 1822 1272 1825 1278
rect 2190 1272 2193 1278
rect 2206 1272 2209 1278
rect 2406 1272 2409 1278
rect 246 1268 398 1271
rect 454 1268 486 1271
rect 490 1268 518 1271
rect 538 1268 622 1271
rect 634 1268 638 1271
rect 650 1268 654 1271
rect 666 1268 670 1271
rect 734 1268 830 1271
rect 890 1268 934 1271
rect 950 1268 974 1271
rect 986 1268 1046 1271
rect 1074 1268 1190 1271
rect 1194 1268 1270 1271
rect 1282 1268 1302 1271
rect 1314 1268 1326 1271
rect 1338 1268 1342 1271
rect 1354 1268 1374 1271
rect 1466 1268 1470 1271
rect 1482 1268 1494 1271
rect 1570 1268 1598 1271
rect 1634 1268 1654 1271
rect 1714 1268 1758 1271
rect 1906 1268 1958 1271
rect 2018 1268 2030 1271
rect 2058 1268 2070 1271
rect 2422 1271 2425 1278
rect 3422 1272 3425 1278
rect 2422 1268 2430 1271
rect 2610 1268 2702 1271
rect 2738 1268 2766 1271
rect 2786 1268 2798 1271
rect 2802 1268 2838 1271
rect 2906 1268 3006 1271
rect 3058 1268 3182 1271
rect 3226 1268 3278 1271
rect 3282 1268 3350 1271
rect 3354 1268 3366 1271
rect 3378 1268 3406 1271
rect 3434 1268 3438 1271
rect 3614 1271 3617 1278
rect 3602 1268 3617 1271
rect 3622 1272 3625 1278
rect 3674 1268 3750 1271
rect 3794 1268 3822 1271
rect 4002 1268 4022 1271
rect 4218 1268 4222 1271
rect 4258 1268 4270 1271
rect 4338 1268 4350 1271
rect 110 1262 113 1268
rect 246 1262 249 1268
rect 454 1262 457 1268
rect 526 1262 529 1268
rect 734 1262 737 1268
rect 162 1258 190 1261
rect 434 1258 454 1261
rect 498 1258 502 1261
rect 570 1258 598 1261
rect 618 1258 678 1261
rect 714 1258 726 1261
rect 830 1261 833 1268
rect 826 1258 833 1261
rect 878 1261 881 1268
rect 842 1258 881 1261
rect 950 1262 953 1268
rect 954 1258 1126 1261
rect 1130 1258 1134 1261
rect 1162 1258 1166 1261
rect 1266 1258 1286 1261
rect 1330 1258 1334 1261
rect 1346 1258 1398 1261
rect 1426 1258 1454 1261
rect 1510 1261 1513 1268
rect 1474 1258 1513 1261
rect 1526 1262 1529 1268
rect 1538 1258 1553 1261
rect 1626 1258 1670 1261
rect 1706 1258 1758 1261
rect 1770 1258 1782 1261
rect 1802 1258 1830 1261
rect 1834 1258 1942 1261
rect 1946 1258 1950 1261
rect 1990 1261 1993 1268
rect 2286 1262 2289 1268
rect 3758 1262 3761 1268
rect 1990 1258 2006 1261
rect 2506 1258 2510 1261
rect 2514 1258 2542 1261
rect 2762 1258 2790 1261
rect 2946 1258 3046 1261
rect 3154 1258 3318 1261
rect 3322 1258 3366 1261
rect 3370 1258 3406 1261
rect 3410 1258 3694 1261
rect 3778 1258 3830 1261
rect 3834 1258 3886 1261
rect 3894 1261 3897 1268
rect 3894 1258 3910 1261
rect 4026 1258 4046 1261
rect 4050 1258 4158 1261
rect 4230 1261 4233 1268
rect 4230 1258 4246 1261
rect 4266 1258 4334 1261
rect 1182 1252 1185 1258
rect 1550 1252 1553 1258
rect -26 1251 -22 1252
rect -26 1248 14 1251
rect 58 1248 110 1251
rect 450 1248 454 1251
rect 458 1248 574 1251
rect 626 1248 630 1251
rect 658 1248 662 1251
rect 682 1248 710 1251
rect 826 1248 846 1251
rect 850 1248 926 1251
rect 954 1248 1081 1251
rect 1098 1248 1182 1251
rect 1210 1248 1358 1251
rect 1402 1248 1422 1251
rect 1490 1248 1494 1251
rect 1506 1248 1542 1251
rect 1618 1248 1630 1251
rect 1642 1248 1910 1251
rect 1986 1248 2062 1251
rect 2094 1248 2590 1251
rect 2594 1248 2998 1251
rect 3074 1248 3118 1251
rect 3162 1248 3254 1251
rect 3314 1248 3334 1251
rect 3354 1248 3382 1251
rect 3402 1248 3510 1251
rect 3522 1248 3542 1251
rect 3586 1248 3646 1251
rect 3650 1248 3718 1251
rect 3722 1248 3846 1251
rect 4014 1251 4017 1258
rect 3874 1248 4017 1251
rect 4022 1252 4025 1258
rect 4042 1248 4046 1251
rect 4126 1248 4134 1251
rect 4358 1251 4361 1258
rect 4330 1248 4361 1251
rect 1078 1242 1081 1248
rect 482 1238 510 1241
rect 514 1238 534 1241
rect 578 1238 798 1241
rect 842 1238 846 1241
rect 1154 1238 1158 1241
rect 1170 1238 1542 1241
rect 1570 1238 1654 1241
rect 1682 1238 1710 1241
rect 2094 1241 2097 1248
rect 1754 1238 2097 1241
rect 2106 1238 2110 1241
rect 2114 1238 2278 1241
rect 2306 1238 2686 1241
rect 2998 1241 3001 1248
rect 2998 1238 3214 1241
rect 3394 1238 3582 1241
rect 3610 1238 3726 1241
rect 3930 1238 3950 1241
rect 4066 1238 4110 1241
rect 4114 1238 4238 1241
rect 4346 1238 4358 1241
rect 366 1231 369 1238
rect 366 1228 582 1231
rect 586 1228 686 1231
rect 746 1228 910 1231
rect 914 1228 1022 1231
rect 1314 1228 1510 1231
rect 1570 1228 1742 1231
rect 1754 1228 1854 1231
rect 1914 1228 1966 1231
rect 2146 1228 2318 1231
rect 2322 1228 2486 1231
rect 2578 1228 3214 1231
rect 3230 1231 3233 1238
rect 3230 1228 3302 1231
rect 3362 1228 3494 1231
rect 3498 1228 3505 1231
rect 3530 1228 3934 1231
rect 4138 1228 4142 1231
rect 458 1218 638 1221
rect 642 1218 918 1221
rect 930 1218 966 1221
rect 970 1218 1102 1221
rect 1106 1218 1110 1221
rect 1146 1218 1166 1221
rect 1250 1218 1606 1221
rect 1626 1218 1662 1221
rect 1770 1218 1862 1221
rect 1914 1218 2054 1221
rect 2138 1218 2254 1221
rect 2258 1218 2558 1221
rect 2610 1218 2622 1221
rect 2626 1218 2710 1221
rect 2978 1218 3014 1221
rect 3018 1218 3102 1221
rect 3106 1218 3950 1221
rect 4114 1218 4174 1221
rect 418 1208 558 1211
rect 618 1208 726 1211
rect 858 1208 870 1211
rect 1042 1208 1134 1211
rect 1162 1208 1406 1211
rect 1498 1208 1606 1211
rect 1610 1208 2350 1211
rect 3098 1208 3126 1211
rect 3242 1208 3398 1211
rect 3402 1208 3446 1211
rect 3530 1208 3822 1211
rect 4034 1208 4062 1211
rect 4066 1208 4078 1211
rect 4082 1208 4238 1211
rect 392 1203 394 1207
rect 398 1203 401 1207
rect 406 1203 408 1207
rect 1416 1203 1418 1207
rect 1422 1203 1425 1207
rect 1430 1203 1432 1207
rect 2440 1203 2442 1207
rect 2446 1203 2449 1207
rect 2454 1203 2456 1207
rect 3472 1203 3474 1207
rect 3478 1203 3481 1207
rect 3486 1203 3488 1207
rect 122 1198 126 1201
rect 418 1198 558 1201
rect 562 1198 566 1201
rect 698 1198 758 1201
rect 770 1198 982 1201
rect 1498 1198 1550 1201
rect 1570 1198 1598 1201
rect 1642 1198 1670 1201
rect 1778 1198 1974 1201
rect 2154 1198 2166 1201
rect 2178 1198 2302 1201
rect 2874 1198 2990 1201
rect 2994 1198 3022 1201
rect 3026 1198 3038 1201
rect 3066 1198 3278 1201
rect 3306 1198 3374 1201
rect 3578 1198 3590 1201
rect 3610 1198 3670 1201
rect 3698 1198 3750 1201
rect 3754 1198 3862 1201
rect 3962 1198 4190 1201
rect 4290 1198 4350 1201
rect 10 1188 798 1191
rect 1310 1191 1313 1198
rect 4198 1192 4201 1198
rect 1310 1188 1334 1191
rect 1338 1188 1494 1191
rect 1514 1188 1662 1191
rect 1666 1188 1742 1191
rect 1818 1188 1894 1191
rect 1898 1188 1918 1191
rect 2098 1188 2102 1191
rect 2106 1188 2198 1191
rect 2594 1188 2910 1191
rect 2930 1188 3174 1191
rect 3226 1188 3238 1191
rect 3242 1188 3294 1191
rect 3298 1188 3406 1191
rect 3410 1188 3566 1191
rect 3586 1188 3654 1191
rect 4022 1188 4030 1191
rect 4034 1188 4182 1191
rect 4242 1188 4382 1191
rect 926 1182 929 1188
rect -26 1181 -22 1182
rect -26 1178 14 1181
rect 378 1178 382 1181
rect 410 1178 454 1181
rect 554 1178 590 1181
rect 706 1178 918 1181
rect 1066 1178 1105 1181
rect 1114 1178 1430 1181
rect 1578 1178 1790 1181
rect 1794 1178 1854 1181
rect 1882 1178 1942 1181
rect 1978 1178 2614 1181
rect 2622 1178 2982 1181
rect 2986 1178 3078 1181
rect 3082 1178 3190 1181
rect 3194 1178 3206 1181
rect 3214 1181 3217 1188
rect 3214 1178 3246 1181
rect 3266 1178 3286 1181
rect 3290 1178 3334 1181
rect 3338 1178 3438 1181
rect 3458 1178 3462 1181
rect 3514 1178 3558 1181
rect 3570 1178 3702 1181
rect 3714 1178 3806 1181
rect 4002 1178 4054 1181
rect 4214 1181 4217 1188
rect 4214 1178 4262 1181
rect 4306 1178 4326 1181
rect 4370 1178 4390 1181
rect 42 1168 94 1171
rect 362 1168 414 1171
rect 434 1168 462 1171
rect 646 1171 649 1178
rect 586 1168 649 1171
rect 754 1168 774 1171
rect 818 1168 1094 1171
rect 1102 1171 1105 1178
rect 1102 1168 1342 1171
rect 1354 1168 1358 1171
rect 1438 1171 1441 1178
rect 2622 1172 2625 1178
rect 1438 1168 1598 1171
rect 1602 1168 1654 1171
rect 1658 1168 1718 1171
rect 1754 1168 1758 1171
rect 1842 1168 1958 1171
rect 2266 1168 2270 1171
rect 2282 1168 2430 1171
rect 2826 1168 2854 1171
rect 2898 1168 2902 1171
rect 3062 1168 3150 1171
rect 3290 1168 3302 1171
rect 3386 1168 3750 1171
rect 3770 1168 3774 1171
rect 3978 1168 4022 1171
rect 4026 1168 4054 1171
rect 4058 1168 4182 1171
rect 4186 1168 4214 1171
rect 4218 1168 4342 1171
rect 4346 1168 4366 1171
rect 422 1161 425 1168
rect 422 1158 502 1161
rect 506 1158 510 1161
rect 566 1161 569 1168
rect 538 1158 638 1161
rect 642 1158 697 1161
rect 706 1158 766 1161
rect 794 1158 854 1161
rect 946 1158 950 1161
rect 1098 1158 1102 1161
rect 1362 1158 1374 1161
rect 1426 1158 1558 1161
rect 1586 1158 1662 1161
rect 1674 1158 1726 1161
rect 1734 1161 1737 1168
rect 1734 1158 1854 1161
rect 1858 1158 1878 1161
rect 1886 1158 1894 1161
rect 1898 1158 1918 1161
rect 1986 1158 2022 1161
rect 2234 1158 2238 1161
rect 2266 1158 2318 1161
rect 2570 1158 2574 1161
rect 2586 1158 2774 1161
rect 2826 1158 2846 1161
rect 2858 1158 2878 1161
rect 2898 1158 2934 1161
rect 3038 1161 3041 1168
rect 3062 1162 3065 1168
rect 3166 1162 3169 1168
rect 3010 1158 3041 1161
rect 3058 1158 3062 1161
rect 3154 1158 3158 1161
rect 3250 1158 3326 1161
rect 3330 1158 3526 1161
rect 3538 1158 3694 1161
rect 3706 1158 3710 1161
rect 3730 1158 3758 1161
rect 3762 1158 3846 1161
rect 3850 1158 3862 1161
rect 3866 1158 3902 1161
rect 3994 1158 3998 1161
rect 4054 1158 4062 1161
rect 4066 1158 4110 1161
rect 4122 1158 4158 1161
rect 4218 1158 4222 1161
rect 4290 1158 4310 1161
rect -26 1151 -22 1152
rect -26 1148 62 1151
rect 86 1151 89 1158
rect 86 1148 134 1151
rect 138 1148 145 1151
rect 162 1148 198 1151
rect 378 1148 438 1151
rect 442 1148 614 1151
rect 682 1148 686 1151
rect 694 1151 697 1158
rect 1062 1152 1065 1158
rect 1070 1152 1073 1158
rect 1118 1152 1121 1158
rect 1126 1152 1129 1158
rect 1142 1152 1145 1158
rect 1326 1152 1329 1158
rect 1334 1152 1337 1158
rect 2214 1152 2217 1158
rect 2814 1152 2817 1158
rect 3046 1152 3049 1158
rect 3102 1152 3105 1158
rect 694 1148 702 1151
rect 722 1148 766 1151
rect 930 1148 950 1151
rect 994 1148 998 1151
rect 1082 1148 1110 1151
rect 1150 1148 1302 1151
rect 1338 1148 1446 1151
rect 1466 1148 1510 1151
rect 1514 1148 1694 1151
rect 1722 1148 1785 1151
rect 1794 1148 1822 1151
rect 1986 1148 1998 1151
rect 2002 1148 2014 1151
rect 2122 1148 2126 1151
rect 2202 1148 2206 1151
rect 2226 1148 2286 1151
rect 2290 1148 2302 1151
rect 2306 1148 2526 1151
rect 2554 1148 2558 1151
rect 2618 1148 2630 1151
rect 2850 1148 2870 1151
rect 2882 1148 2926 1151
rect 2938 1148 3046 1151
rect 3074 1148 3078 1151
rect 3114 1148 3118 1151
rect 3134 1151 3137 1158
rect 3134 1148 3142 1151
rect 3162 1148 3198 1151
rect 3250 1148 3254 1151
rect 3258 1148 3414 1151
rect 3418 1148 3478 1151
rect 3498 1148 3502 1151
rect 3546 1148 3606 1151
rect 3626 1148 3630 1151
rect 3722 1148 3726 1151
rect 3754 1148 3769 1151
rect 3778 1148 3782 1151
rect 3930 1148 4030 1151
rect 4058 1148 4070 1151
rect 4090 1148 4126 1151
rect 4154 1148 4294 1151
rect 4338 1148 4358 1151
rect 806 1142 809 1148
rect 378 1138 534 1141
rect 538 1138 718 1141
rect 850 1138 934 1141
rect 954 1138 982 1141
rect 1150 1141 1153 1148
rect 1002 1138 1153 1141
rect 1214 1138 1230 1141
rect 1282 1138 1382 1141
rect 1466 1138 1470 1141
rect 1490 1138 1510 1141
rect 1514 1138 1718 1141
rect 1782 1141 1785 1148
rect 3678 1142 3681 1148
rect 3766 1142 3769 1148
rect 1782 1138 1846 1141
rect 1850 1138 1862 1141
rect 1882 1138 3190 1141
rect 3194 1138 3398 1141
rect 3402 1138 3478 1141
rect 3482 1138 3614 1141
rect 3798 1141 3801 1148
rect 3798 1138 3822 1141
rect 3826 1138 3926 1141
rect 3938 1138 3958 1141
rect 3962 1138 4006 1141
rect 4010 1138 4038 1141
rect 4042 1138 4166 1141
rect 4170 1138 4198 1141
rect 4202 1138 4326 1141
rect 1214 1132 1217 1138
rect 466 1128 494 1131
rect 498 1128 606 1131
rect 650 1128 654 1131
rect 674 1128 750 1131
rect 786 1128 886 1131
rect 890 1128 1086 1131
rect 1106 1128 1206 1131
rect 1298 1128 1489 1131
rect 1498 1128 1502 1131
rect 1530 1128 1534 1131
rect 1546 1128 1550 1131
rect 1570 1128 1630 1131
rect 1634 1128 1718 1131
rect 1818 1128 1822 1131
rect 1834 1128 1862 1131
rect 1866 1128 1870 1131
rect 1954 1128 1958 1131
rect 2002 1128 2006 1131
rect 2018 1128 2198 1131
rect 2206 1128 2222 1131
rect 2238 1128 2286 1131
rect 2314 1128 2342 1131
rect 2346 1128 2398 1131
rect 2530 1128 2574 1131
rect 2586 1128 2614 1131
rect 2718 1128 2814 1131
rect 2818 1128 2990 1131
rect 3082 1128 3086 1131
rect 3098 1128 3150 1131
rect 3202 1128 3206 1131
rect 3226 1128 3230 1131
rect 3238 1128 3278 1131
rect 3322 1128 3350 1131
rect 3378 1128 3414 1131
rect 3418 1128 3462 1131
rect 3506 1128 3694 1131
rect 3758 1131 3761 1138
rect 3722 1128 3761 1131
rect 3818 1128 3838 1131
rect 3882 1128 3886 1131
rect 4098 1128 4190 1131
rect 4306 1128 4326 1131
rect 270 1122 273 1128
rect 1230 1122 1233 1128
rect 130 1118 222 1121
rect 298 1118 382 1121
rect 426 1118 542 1121
rect 578 1118 678 1121
rect 710 1118 718 1121
rect 722 1118 798 1121
rect 906 1118 934 1121
rect 954 1118 1046 1121
rect 1058 1118 1206 1121
rect 1250 1118 1350 1121
rect 1354 1118 1374 1121
rect 1402 1118 1478 1121
rect 1486 1121 1489 1128
rect 1590 1122 1593 1128
rect 1486 1118 1502 1121
rect 1514 1118 1582 1121
rect 1610 1118 1622 1121
rect 1650 1118 1654 1121
rect 1674 1118 1678 1121
rect 1698 1118 1710 1121
rect 1750 1121 1753 1128
rect 1750 1118 1902 1121
rect 1906 1118 1918 1121
rect 2006 1121 2009 1128
rect 2206 1122 2209 1128
rect 2238 1122 2241 1128
rect 2718 1122 2721 1128
rect 2006 1118 2014 1121
rect 2106 1118 2134 1121
rect 2154 1118 2190 1121
rect 2250 1118 2254 1121
rect 2322 1118 2390 1121
rect 2450 1118 2654 1121
rect 2738 1118 2742 1121
rect 2834 1118 2846 1121
rect 2930 1118 2950 1121
rect 2954 1118 2998 1121
rect 3006 1118 3009 1128
rect 3158 1121 3161 1128
rect 3018 1118 3161 1121
rect 3238 1122 3241 1128
rect 4070 1122 4073 1128
rect 4270 1122 4273 1128
rect 3250 1118 3286 1121
rect 3298 1118 3390 1121
rect 3522 1118 3526 1121
rect 3698 1118 3886 1121
rect 4090 1118 4158 1121
rect 2862 1112 2865 1118
rect 154 1108 614 1111
rect 970 1108 1022 1111
rect 1026 1108 1110 1111
rect 1114 1108 1166 1111
rect 1258 1108 1262 1111
rect 1322 1108 1350 1111
rect 1362 1108 1374 1111
rect 1386 1108 1390 1111
rect 1426 1108 1822 1111
rect 2026 1108 2166 1111
rect 2202 1108 2350 1111
rect 2394 1108 2398 1111
rect 2426 1108 2438 1111
rect 2586 1108 2766 1111
rect 2898 1108 2942 1111
rect 2986 1108 3118 1111
rect 3122 1108 3350 1111
rect 3402 1108 3422 1111
rect 3426 1108 3462 1111
rect 3562 1108 3622 1111
rect 3714 1108 3718 1111
rect 3730 1108 3942 1111
rect 4266 1108 4366 1111
rect 734 1102 737 1108
rect 862 1102 865 1108
rect 896 1103 898 1107
rect 902 1103 905 1107
rect 910 1103 912 1107
rect 1928 1103 1930 1107
rect 1934 1103 1937 1107
rect 1942 1103 1944 1107
rect 186 1098 190 1101
rect 258 1098 550 1101
rect 674 1098 678 1101
rect 946 1098 1430 1101
rect 1466 1098 1470 1101
rect 1474 1098 1486 1101
rect 1522 1098 1550 1101
rect 1554 1098 1614 1101
rect 1618 1098 1702 1101
rect 1706 1098 1734 1101
rect 1850 1098 1878 1101
rect 1954 1098 2094 1101
rect 2098 1098 2118 1101
rect 2298 1098 2342 1101
rect 2350 1101 2353 1108
rect 2952 1103 2954 1107
rect 2958 1103 2961 1107
rect 2966 1103 2968 1107
rect 3976 1103 3978 1107
rect 3982 1103 3985 1107
rect 3990 1103 3992 1107
rect 2350 1098 2534 1101
rect 2546 1098 2830 1101
rect 2834 1098 2926 1101
rect 2994 1098 3134 1101
rect 3146 1098 3198 1101
rect 3250 1098 3550 1101
rect 3658 1098 3742 1101
rect 3998 1098 4198 1101
rect 4258 1098 4294 1101
rect 4346 1098 4358 1101
rect 282 1088 366 1091
rect 538 1088 854 1091
rect 874 1088 1001 1091
rect 1010 1088 1334 1091
rect 1354 1088 1406 1091
rect 1450 1088 1510 1091
rect 1530 1088 1534 1091
rect 1538 1088 1550 1091
rect 1566 1088 1574 1091
rect 1578 1088 1630 1091
rect 1642 1088 1774 1091
rect 1778 1088 1870 1091
rect 1874 1088 1894 1091
rect 1898 1088 1918 1091
rect 1922 1088 2382 1091
rect 2402 1088 2606 1091
rect 2610 1088 2638 1091
rect 2706 1088 3518 1091
rect 3522 1088 3542 1091
rect 3714 1088 3766 1091
rect 3998 1091 4001 1098
rect 3986 1088 4001 1091
rect 4178 1088 4206 1091
rect 4314 1088 4358 1091
rect 6 1081 9 1088
rect 998 1082 1001 1088
rect 2062 1082 2065 1088
rect 2462 1082 2465 1088
rect 3622 1082 3625 1088
rect -26 1078 9 1081
rect 370 1078 430 1081
rect 442 1078 518 1081
rect 546 1078 654 1081
rect 666 1078 766 1081
rect 802 1078 950 1081
rect 1274 1078 1278 1081
rect 1330 1078 1345 1081
rect 1370 1078 1566 1081
rect 1578 1078 1582 1081
rect 1626 1078 1646 1081
rect 1690 1078 1710 1081
rect 1806 1078 1814 1081
rect 1818 1078 1822 1081
rect 1854 1078 1862 1081
rect 1902 1078 1910 1081
rect 1914 1078 1966 1081
rect 1978 1078 1982 1081
rect 2026 1078 2030 1081
rect 2122 1078 2126 1081
rect 2170 1078 2222 1081
rect 2254 1078 2318 1081
rect 2330 1078 2430 1081
rect 2538 1078 2542 1081
rect 2546 1078 2590 1081
rect 2602 1078 2654 1081
rect 2682 1078 2718 1081
rect 2758 1078 2774 1081
rect 2866 1078 2886 1081
rect 2890 1078 2894 1081
rect 2938 1078 2958 1081
rect 3146 1078 3206 1081
rect 3210 1078 3214 1081
rect 3218 1078 3278 1081
rect 3290 1078 3342 1081
rect 3458 1078 3470 1081
rect 3514 1078 3566 1081
rect 3578 1078 3582 1081
rect 3674 1078 3694 1081
rect 3702 1081 3705 1088
rect 3702 1078 3726 1081
rect 3730 1078 3742 1081
rect 3838 1081 3841 1088
rect 3838 1078 3902 1081
rect 3906 1078 3942 1081
rect 4138 1078 4190 1081
rect 4202 1078 4302 1081
rect 4378 1078 4390 1081
rect -26 1072 -23 1078
rect -26 1068 -22 1072
rect 30 1071 33 1078
rect 10 1068 33 1071
rect 142 1072 145 1078
rect 158 1072 161 1078
rect 1070 1072 1073 1078
rect 610 1068 638 1071
rect 658 1068 726 1071
rect 730 1068 734 1071
rect 770 1068 990 1071
rect 1002 1068 1014 1071
rect 1274 1068 1278 1071
rect 1342 1071 1345 1078
rect 1342 1068 1385 1071
rect 414 1062 417 1068
rect 1046 1062 1049 1068
rect 34 1058 246 1061
rect 426 1058 462 1061
rect 650 1058 662 1061
rect 746 1058 750 1061
rect 906 1058 966 1061
rect 986 1058 990 1061
rect 1010 1058 1046 1061
rect 1178 1058 1294 1061
rect 1302 1061 1305 1068
rect 1334 1061 1337 1068
rect 1302 1058 1337 1061
rect 1382 1062 1385 1068
rect 1470 1068 1478 1071
rect 1482 1068 1526 1071
rect 1538 1068 1542 1071
rect 1766 1071 1769 1078
rect 1854 1072 1857 1078
rect 1554 1068 1769 1071
rect 1778 1068 1790 1071
rect 1810 1068 1814 1071
rect 1866 1068 1926 1071
rect 1954 1068 2078 1071
rect 2254 1071 2257 1078
rect 2758 1072 2761 1078
rect 2106 1068 2257 1071
rect 2266 1068 2406 1071
rect 2410 1068 2478 1071
rect 2546 1068 2550 1071
rect 2554 1068 2670 1071
rect 2706 1068 2758 1071
rect 2826 1068 2870 1071
rect 2918 1071 2921 1078
rect 3094 1072 3097 1078
rect 3110 1072 3113 1078
rect 2918 1068 2934 1071
rect 2946 1068 2974 1071
rect 3186 1068 3310 1071
rect 3338 1068 3366 1071
rect 3370 1068 3414 1071
rect 3438 1071 3441 1078
rect 3790 1072 3793 1078
rect 4134 1072 4137 1078
rect 4342 1072 4345 1078
rect 3418 1068 3441 1071
rect 3450 1068 3574 1071
rect 3634 1068 3654 1071
rect 3690 1068 3718 1071
rect 3738 1068 3742 1071
rect 3946 1068 3958 1071
rect 3978 1068 4102 1071
rect 4154 1068 4166 1071
rect 4194 1068 4198 1071
rect 4242 1068 4310 1071
rect 1406 1062 1409 1068
rect 1438 1061 1441 1068
rect 3598 1062 3601 1068
rect 1438 1058 1462 1061
rect 1482 1058 1486 1061
rect 1514 1058 1566 1061
rect 1586 1058 1638 1061
rect 1666 1058 1686 1061
rect 1730 1058 1950 1061
rect 2058 1058 2094 1061
rect 2142 1058 2390 1061
rect 2562 1058 2622 1061
rect 2658 1058 2774 1061
rect 2938 1058 2942 1061
rect 2978 1058 3006 1061
rect 3010 1058 3198 1061
rect 3250 1058 3262 1061
rect 3266 1058 3342 1061
rect 3346 1058 3374 1061
rect 3378 1058 3446 1061
rect 3514 1058 3542 1061
rect 3570 1058 3574 1061
rect 3650 1058 3662 1061
rect 3682 1058 3790 1061
rect 3946 1058 3966 1061
rect 4066 1058 4094 1061
rect 4146 1058 4150 1061
rect 4162 1058 4166 1061
rect 4186 1058 4270 1061
rect 4290 1058 4326 1061
rect 1078 1052 1081 1058
rect 1646 1052 1649 1058
rect 2142 1052 2145 1058
rect 2478 1052 2481 1058
rect 3470 1052 3473 1058
rect -26 1051 -22 1052
rect -26 1048 6 1051
rect 354 1048 430 1051
rect 522 1048 662 1051
rect 682 1048 702 1051
rect 722 1048 753 1051
rect 770 1048 774 1051
rect 866 1048 1054 1051
rect 1154 1048 1278 1051
rect 1306 1048 1350 1051
rect 1394 1048 1582 1051
rect 1594 1048 1606 1051
rect 1682 1048 1686 1051
rect 1826 1048 1830 1051
rect 1834 1048 1854 1051
rect 1858 1048 2030 1051
rect 2034 1048 2094 1051
rect 2282 1048 2286 1051
rect 2322 1048 2350 1051
rect 2370 1048 2374 1051
rect 2666 1048 2686 1051
rect 2866 1048 2958 1051
rect 3226 1048 3358 1051
rect 3362 1048 3374 1051
rect 3482 1048 3502 1051
rect 3602 1048 3702 1051
rect 4018 1048 4022 1051
rect 4026 1048 4046 1051
rect 4050 1048 4078 1051
rect 4082 1048 4158 1051
rect 4162 1048 4238 1051
rect 4274 1048 4294 1051
rect 4298 1048 4302 1051
rect 750 1042 753 1048
rect 1806 1042 1809 1048
rect 3598 1042 3601 1048
rect 666 1038 670 1041
rect 706 1038 726 1041
rect 822 1038 1174 1041
rect 1314 1038 1542 1041
rect 1570 1038 1638 1041
rect 1874 1038 1990 1041
rect 1994 1038 2382 1041
rect 2386 1038 2422 1041
rect 2434 1038 3238 1041
rect 3354 1038 3558 1041
rect 3650 1038 3702 1041
rect 3966 1041 3969 1048
rect 3966 1038 3998 1041
rect 4034 1038 4062 1041
rect 4066 1038 4094 1041
rect 4098 1038 4134 1041
rect 4138 1038 4238 1041
rect 4242 1038 4246 1041
rect 822 1031 825 1038
rect 4270 1032 4273 1038
rect 434 1028 825 1031
rect 922 1028 1054 1031
rect 1146 1028 1590 1031
rect 1602 1028 1782 1031
rect 1890 1028 3006 1031
rect 3010 1028 3494 1031
rect 3578 1028 3662 1031
rect 3826 1028 4006 1031
rect 4098 1028 4102 1031
rect 4154 1028 4174 1031
rect 4226 1028 4230 1031
rect 674 1018 710 1021
rect 714 1018 721 1021
rect 1034 1018 1038 1021
rect 1066 1018 1441 1021
rect 1466 1018 1470 1021
rect 1586 1018 1758 1021
rect 1762 1018 1942 1021
rect 1954 1018 2006 1021
rect 2130 1018 2246 1021
rect 2326 1018 2486 1021
rect 2490 1018 4070 1021
rect 4210 1018 4222 1021
rect 530 1008 534 1011
rect 690 1008 878 1011
rect 882 1008 886 1011
rect 1018 1008 1038 1011
rect 1058 1008 1070 1011
rect 1170 1008 1374 1011
rect 1378 1008 1390 1011
rect 1438 1011 1441 1018
rect 1574 1012 1577 1018
rect 2326 1012 2329 1018
rect 1438 1008 1534 1011
rect 1818 1008 1862 1011
rect 1882 1008 1910 1011
rect 1962 1008 2046 1011
rect 2146 1008 2214 1011
rect 2218 1008 2326 1011
rect 2346 1008 2358 1011
rect 2738 1008 3022 1011
rect 3090 1008 3110 1011
rect 3290 1008 3342 1011
rect 3346 1008 3390 1011
rect 3578 1008 3622 1011
rect 3842 1008 4038 1011
rect 392 1003 394 1007
rect 398 1003 401 1007
rect 406 1003 408 1007
rect 1416 1003 1418 1007
rect 1422 1003 1425 1007
rect 1430 1003 1432 1007
rect 2440 1003 2442 1007
rect 2446 1003 2449 1007
rect 2454 1003 2456 1007
rect 3472 1003 3474 1007
rect 3478 1003 3481 1007
rect 3486 1003 3488 1007
rect 4070 1002 4073 1008
rect 1002 998 1094 1001
rect 1138 998 1142 1001
rect 1178 998 1374 1001
rect 1586 998 1694 1001
rect 1922 998 2366 1001
rect 2522 998 2670 1001
rect 2674 998 3014 1001
rect 3114 998 3369 1001
rect -26 991 -22 992
rect -26 988 38 991
rect 298 988 302 991
rect 786 988 1046 991
rect 1050 988 1214 991
rect 1218 988 1654 991
rect 1698 988 1790 991
rect 1994 988 2593 991
rect 2602 988 2606 991
rect 2642 988 2854 991
rect 3242 988 3270 991
rect 3366 991 3369 998
rect 3826 998 3854 1001
rect 3718 992 3721 998
rect 3366 988 3534 991
rect 3562 988 3630 991
rect 3738 988 3798 991
rect 3802 988 3966 991
rect 3970 988 4086 991
rect 262 981 265 988
rect 18 978 265 981
rect 394 978 478 981
rect 730 978 1022 981
rect 1026 978 1030 981
rect 1042 978 1198 981
rect 1322 978 1342 981
rect 1346 978 1574 981
rect 1722 978 1774 981
rect 1786 978 1998 981
rect 2042 978 2102 981
rect 2106 978 2142 981
rect 2242 978 2358 981
rect 2434 978 2542 981
rect 2590 981 2593 988
rect 2894 982 2897 988
rect 2590 978 2742 981
rect 2746 978 2758 981
rect 3158 981 3161 988
rect 3158 978 3438 981
rect 3442 978 3614 981
rect 3618 978 4022 981
rect -26 971 -22 972
rect 6 971 9 978
rect -26 968 9 971
rect 290 968 478 971
rect 1022 968 1166 971
rect 1346 968 2134 971
rect 2138 968 2182 971
rect 2186 968 2390 971
rect 2754 968 2790 971
rect 2794 968 2926 971
rect 2930 968 3118 971
rect 3170 968 3294 971
rect 3458 968 3518 971
rect 3530 968 3710 971
rect 3722 968 3854 971
rect 3874 968 3926 971
rect 4058 968 4094 971
rect 4242 968 4246 971
rect 238 961 241 968
rect 1022 962 1025 968
rect 1326 962 1329 968
rect 26 958 241 961
rect 266 958 294 961
rect 874 958 894 961
rect 1106 958 1110 961
rect 1442 958 1446 961
rect 1450 958 1478 961
rect 1506 958 1510 961
rect 1538 958 1558 961
rect 1642 958 1670 961
rect 1730 958 1742 961
rect 1778 958 1846 961
rect 1850 958 1878 961
rect 1986 958 2022 961
rect 2050 958 2054 961
rect 2478 961 2481 968
rect 2478 958 2502 961
rect 2622 961 2625 968
rect 2554 958 2625 961
rect 2634 958 2734 961
rect 2874 958 2894 961
rect 2898 958 2918 961
rect 3090 958 3238 961
rect 3322 958 3510 961
rect 3518 958 3598 961
rect 3626 958 3782 961
rect 3786 958 3878 961
rect 3962 958 3993 961
rect 4098 958 4198 961
rect 4210 958 4214 961
rect 4250 958 4254 961
rect 1182 952 1185 958
rect -26 951 -22 952
rect -26 948 14 951
rect 162 948 542 951
rect 622 948 742 951
rect 978 948 1006 951
rect 1058 948 1065 951
rect 1074 948 1126 951
rect 1130 948 1142 951
rect 1154 948 1158 951
rect 1198 951 1201 958
rect 1206 951 1209 958
rect 1198 948 1209 951
rect 1222 952 1225 958
rect 1286 952 1289 958
rect 1350 952 1353 958
rect 1250 948 1254 951
rect 1266 948 1270 951
rect 1298 948 1350 951
rect 1358 951 1361 958
rect 1758 952 1761 958
rect 1358 948 1366 951
rect 1378 948 1486 951
rect 1586 948 1702 951
rect 1794 948 1798 951
rect 1858 948 1870 951
rect 1874 948 1878 951
rect 1882 948 1894 951
rect 1898 948 1926 951
rect 1982 951 1985 958
rect 1970 948 1985 951
rect 2042 948 2078 951
rect 2114 948 2118 951
rect 2358 951 2361 958
rect 2358 948 2470 951
rect 2506 948 2510 951
rect 2634 948 2662 951
rect 2770 948 2774 951
rect 2810 948 2814 951
rect 2850 948 3118 951
rect 3130 948 3134 951
rect 442 938 510 941
rect 514 938 526 941
rect 582 941 585 948
rect 622 942 625 948
rect 582 938 590 941
rect 642 938 662 941
rect 806 941 809 948
rect 1006 942 1009 948
rect 706 938 809 941
rect 858 938 902 941
rect 1050 938 1062 941
rect 1090 938 1094 941
rect 1130 938 1134 941
rect 1146 938 1222 941
rect 1230 941 1233 948
rect 1226 938 1233 941
rect 1242 938 1430 941
rect 1434 938 1446 941
rect 1450 938 1478 941
rect 1490 938 1494 941
rect 1570 938 1598 941
rect 1762 938 1790 941
rect 1826 938 1830 941
rect 1858 938 2014 941
rect 2066 938 2150 941
rect 2162 938 2166 941
rect 2170 938 2198 941
rect 2346 938 2366 941
rect 2370 938 2406 941
rect 2410 938 2470 941
rect 2474 938 2510 941
rect 2534 941 2537 948
rect 2750 942 2753 948
rect 2530 938 2537 941
rect 2626 938 2678 941
rect 2690 938 2734 941
rect 2890 938 3134 941
rect 3146 938 3150 941
rect 3198 941 3201 948
rect 3154 938 3201 941
rect 3394 948 3398 951
rect 3422 948 3462 951
rect 3518 951 3521 958
rect 3990 952 3993 958
rect 3482 948 3521 951
rect 3586 948 3622 951
rect 3658 948 3662 951
rect 3762 948 3766 951
rect 3842 948 3926 951
rect 3998 948 4030 951
rect 4046 948 4062 951
rect 4114 948 4118 951
rect 4170 948 4182 951
rect 4234 948 4254 951
rect 3294 941 3297 948
rect 3422 942 3425 948
rect 3774 942 3777 948
rect 3998 942 4001 948
rect 4046 942 4049 948
rect 3294 938 3350 941
rect 3458 938 3542 941
rect 3546 938 3734 941
rect 3742 938 3750 941
rect 3818 938 3822 941
rect 3922 938 3950 941
rect 4058 938 4094 941
rect 4122 938 4126 941
rect 4130 938 4222 941
rect 4250 938 4254 941
rect 4266 938 4270 941
rect 4290 938 4358 941
rect 142 928 150 931
rect 658 928 713 931
rect 778 928 793 931
rect 1010 928 1070 931
rect 1098 928 1150 931
rect 1154 928 1262 931
rect 1266 928 1294 931
rect 1346 928 1382 931
rect 1510 931 1513 938
rect 1482 928 1513 931
rect 1530 928 1606 931
rect 1642 928 1646 931
rect 1742 931 1745 938
rect 2678 932 2681 938
rect 3414 932 3417 938
rect 1706 928 1745 931
rect 1762 928 1806 931
rect 1858 928 1878 931
rect 1922 928 1926 931
rect 1946 928 2118 931
rect 2130 928 2134 931
rect 2138 928 2150 931
rect 2258 928 2350 931
rect 2402 928 2422 931
rect 2450 928 2494 931
rect 2502 928 2598 931
rect 2834 928 2846 931
rect 2874 928 2910 931
rect 3130 928 3294 931
rect 3314 928 3326 931
rect 3330 928 3366 931
rect 3426 928 3462 931
rect 3522 928 3550 931
rect 3554 928 3710 931
rect 3714 928 3806 931
rect 3818 928 3910 931
rect 4010 928 4022 931
rect 4026 928 4038 931
rect 4042 928 4086 931
rect 4090 928 4198 931
rect 4202 928 4222 931
rect 4274 928 4326 931
rect 142 922 145 928
rect 374 922 377 928
rect 710 922 713 928
rect 790 922 793 928
rect 850 918 1022 921
rect 1042 918 1166 921
rect 1218 918 1230 921
rect 1266 918 1342 921
rect 1362 918 1366 921
rect 1466 918 1558 921
rect 1578 918 1614 921
rect 1642 918 1742 921
rect 1746 918 1958 921
rect 1978 918 1982 921
rect 1994 918 2094 921
rect 2374 921 2377 928
rect 2374 918 2382 921
rect 2502 921 2505 928
rect 2418 918 2505 921
rect 2514 918 2534 921
rect 2538 918 2590 921
rect 2594 918 2646 921
rect 2650 918 2710 921
rect 2810 918 2902 921
rect 2922 918 2942 921
rect 3050 918 3198 921
rect 3378 918 3446 921
rect 3450 918 3590 921
rect 3610 918 3622 921
rect 3626 918 3633 921
rect 3642 918 3694 921
rect 3698 918 3710 921
rect 3714 918 3742 921
rect 3762 918 3790 921
rect 3914 918 3942 921
rect 3986 918 3998 921
rect 4010 918 4182 921
rect 4186 918 4198 921
rect 4262 918 4286 921
rect 682 908 710 911
rect 794 908 886 911
rect 946 908 1086 911
rect 1122 908 1126 911
rect 1290 908 1454 911
rect 1498 908 1502 911
rect 1522 908 1550 911
rect 1586 908 1886 911
rect 1994 908 2238 911
rect 2378 908 2390 911
rect 2458 908 2502 911
rect 2506 908 2614 911
rect 2682 908 2806 911
rect 2818 908 2830 911
rect 3090 908 3102 911
rect 3130 908 3262 911
rect 3290 908 3382 911
rect 3386 908 3406 911
rect 3410 908 3414 911
rect 3638 911 3641 918
rect 3418 908 3641 911
rect 3650 908 3790 911
rect 4002 908 4070 911
rect 4262 911 4265 918
rect 4186 908 4265 911
rect 4274 908 4278 911
rect 896 903 898 907
rect 902 903 905 907
rect 910 903 912 907
rect 1928 903 1930 907
rect 1934 903 1937 907
rect 1942 903 1944 907
rect 2952 903 2954 907
rect 2958 903 2961 907
rect 2966 903 2968 907
rect 3976 903 3978 907
rect 3982 903 3985 907
rect 3990 903 3992 907
rect 570 898 766 901
rect 778 898 854 901
rect 922 898 1318 901
rect 1330 898 1334 901
rect 1394 898 1526 901
rect 1530 898 1558 901
rect 1562 898 1614 901
rect 1690 898 1718 901
rect 2050 898 2310 901
rect 2354 898 2566 901
rect 2594 898 2614 901
rect 2826 898 2838 901
rect 2842 898 2926 901
rect 2930 898 2942 901
rect 3058 898 3230 901
rect 3266 898 3278 901
rect 3282 898 3526 901
rect 3746 898 3846 901
rect 4066 898 4078 901
rect 4082 898 4126 901
rect 4130 898 4158 901
rect 4258 898 4318 901
rect 614 888 622 891
rect 626 888 774 891
rect 778 888 1110 891
rect 1114 888 1134 891
rect 1306 888 1326 891
rect 1330 888 1337 891
rect 1346 888 1390 891
rect 1458 888 1462 891
rect 1474 888 1502 891
rect 1546 888 1582 891
rect 1722 888 1726 891
rect 2002 888 2481 891
rect 2490 888 2601 891
rect 2610 888 2878 891
rect 2882 888 2966 891
rect 2970 888 3046 891
rect 3050 888 3094 891
rect 3122 888 3126 891
rect 3146 888 3174 891
rect 3178 888 3182 891
rect 3314 888 3438 891
rect 3538 888 3542 891
rect 3554 888 3622 891
rect 3626 888 3718 891
rect 3726 888 3798 891
rect 3866 888 4006 891
rect 4194 888 4257 891
rect 142 881 145 888
rect 142 878 262 881
rect 266 878 422 881
rect 458 878 678 881
rect 722 878 758 881
rect 794 878 798 881
rect 818 878 982 881
rect 994 878 1014 881
rect 1154 878 1286 881
rect 1298 878 1310 881
rect 1314 878 1350 881
rect 1406 881 1409 888
rect 1406 878 1510 881
rect 1514 878 1542 881
rect 1626 878 1646 881
rect 1702 881 1705 888
rect 1702 878 1718 881
rect 1762 878 1782 881
rect 1802 878 1806 881
rect 1826 878 1830 881
rect 1850 878 1886 881
rect 1982 881 1985 888
rect 2478 882 2481 888
rect 2598 882 2601 888
rect 1890 878 1985 881
rect 2090 878 2094 881
rect 2378 878 2430 881
rect 2498 878 2518 881
rect 2530 878 2582 881
rect 2586 878 2590 881
rect 2618 878 2622 881
rect 2666 878 2670 881
rect 2698 878 2785 881
rect -26 871 -22 872
rect 6 871 9 878
rect 1734 872 1737 878
rect 2222 872 2225 878
rect 2782 872 2785 878
rect 2842 878 2873 881
rect 2946 878 2974 881
rect 3110 881 3113 888
rect 3726 882 3729 888
rect 4254 882 4257 888
rect 3082 878 3113 881
rect 3118 878 3225 881
rect -26 868 9 871
rect 242 868 302 871
rect 378 868 550 871
rect 690 868 734 871
rect 770 868 926 871
rect 1018 868 1022 871
rect 1146 868 1358 871
rect 1466 868 1510 871
rect 1546 868 1574 871
rect 1578 868 1638 871
rect 1682 868 1686 871
rect 1714 868 1718 871
rect 1770 868 1774 871
rect 1794 868 1814 871
rect 1818 868 1846 871
rect 1978 868 1982 871
rect 2058 868 2166 871
rect 2314 868 2350 871
rect 2402 868 2406 871
rect 2426 868 2574 871
rect 2578 868 2590 871
rect 2594 868 2662 871
rect 2666 868 2750 871
rect 2794 868 2798 871
rect 2822 871 2825 878
rect 2870 872 2873 878
rect 2822 868 2854 871
rect 2898 868 2982 871
rect 2986 868 3006 871
rect 3118 871 3121 878
rect 3222 872 3225 878
rect 3346 878 3374 881
rect 3434 878 3662 881
rect 3706 878 3718 881
rect 3738 878 3782 881
rect 3826 878 3862 881
rect 3946 878 4022 881
rect 4122 878 4150 881
rect 4170 878 4174 881
rect 4190 878 4198 881
rect 4322 878 4350 881
rect 3246 872 3249 878
rect 3098 868 3121 871
rect 3138 868 3182 871
rect 3422 871 3425 878
rect 3358 868 3425 871
rect 3434 868 3462 871
rect 3482 868 3742 871
rect 3770 868 3806 871
rect 3850 868 3934 871
rect 3938 868 4014 871
rect 4018 868 4030 871
rect 4094 871 4097 878
rect 4190 872 4193 878
rect 4094 868 4118 871
rect 4130 868 4134 871
rect 158 862 161 868
rect -26 858 30 861
rect 258 858 654 861
rect 686 861 689 868
rect 2766 862 2769 868
rect 3334 862 3337 868
rect 682 858 689 861
rect 754 858 758 861
rect 762 858 806 861
rect 826 858 830 861
rect 914 858 1038 861
rect 1314 858 1318 861
rect 1322 858 1366 861
rect 1466 858 1478 861
rect 1482 858 1662 861
rect 1666 858 1694 861
rect 1698 858 1702 861
rect 1730 858 1894 861
rect 1898 858 2294 861
rect 2410 858 2414 861
rect 2442 858 2486 861
rect 2522 858 2550 861
rect 2626 858 2630 861
rect 2794 858 2806 861
rect 2874 858 2894 861
rect 2898 858 2990 861
rect 2994 858 3158 861
rect 3242 858 3246 861
rect 3358 861 3361 868
rect 3346 858 3361 861
rect 3370 858 3390 861
rect 3402 858 3406 861
rect 3514 858 3702 861
rect 3714 858 3782 861
rect 3818 858 3830 861
rect 3898 858 3902 861
rect 3914 858 3998 861
rect 4014 861 4017 868
rect 4078 861 4081 868
rect 4206 862 4209 868
rect 4310 862 4313 868
rect 4014 858 4190 861
rect 4234 858 4246 861
rect 4250 858 4286 861
rect -26 852 -23 858
rect -26 848 -22 852
rect 26 848 54 851
rect 522 848 550 851
rect 562 848 753 851
rect 762 848 974 851
rect 1042 848 1366 851
rect 1386 848 1390 851
rect 1394 848 1750 851
rect 1754 848 1870 851
rect 1938 848 1942 851
rect 2302 851 2305 858
rect 2654 852 2657 858
rect 2302 848 2462 851
rect 2466 848 2558 851
rect 2562 848 2622 851
rect 2666 848 2806 851
rect 2810 848 2886 851
rect 2898 848 2902 851
rect 2922 848 2926 851
rect 2938 848 2950 851
rect 3042 848 3070 851
rect 3234 848 3238 851
rect 3266 848 3518 851
rect 3586 848 3766 851
rect 3782 851 3785 858
rect 3782 848 3870 851
rect 3930 848 3934 851
rect 3962 848 3974 851
rect 4018 848 4142 851
rect 4154 848 4166 851
rect 4242 848 4270 851
rect 4282 848 4286 851
rect 4302 851 4305 858
rect 4302 848 4326 851
rect 4330 848 4334 851
rect 238 841 241 848
rect 50 838 241 841
rect 330 838 366 841
rect 370 838 694 841
rect 706 838 718 841
rect 750 841 753 848
rect 3022 842 3025 848
rect 4366 842 4369 848
rect 750 838 966 841
rect 978 838 1310 841
rect 1378 838 1454 841
rect 1498 838 1510 841
rect 1586 838 1590 841
rect 1598 838 1654 841
rect 1666 838 1670 841
rect 1706 838 1710 841
rect 1794 838 1798 841
rect 1810 838 1822 841
rect 1938 838 2046 841
rect 2050 838 2070 841
rect 2090 838 2342 841
rect 2370 838 2494 841
rect 2578 838 2782 841
rect 2786 838 2974 841
rect 3074 838 3174 841
rect 3178 838 3190 841
rect 3202 838 3278 841
rect 3282 838 3286 841
rect 3498 838 3502 841
rect 3898 838 3918 841
rect 4010 838 4038 841
rect 4138 838 4294 841
rect 4334 838 4342 841
rect 694 831 697 838
rect 1598 832 1601 838
rect 2566 832 2569 838
rect 694 828 1030 831
rect 1226 828 1366 831
rect 1674 828 1782 831
rect 1810 828 1862 831
rect 1906 828 1910 831
rect 2370 828 2462 831
rect 2634 828 2774 831
rect 2906 828 3054 831
rect 3082 828 3089 831
rect 3170 828 3174 831
rect 3358 831 3361 838
rect 3218 828 3361 831
rect 3470 831 3473 838
rect 4334 832 4337 838
rect 3426 828 3473 831
rect 3754 828 3806 831
rect 3866 828 3966 831
rect 4042 828 4110 831
rect 4154 828 4326 831
rect 690 818 726 821
rect 930 818 1118 821
rect 1122 818 1270 821
rect 1274 818 1398 821
rect 1434 818 2286 821
rect 2314 818 2414 821
rect 2418 818 2454 821
rect 2602 818 2622 821
rect 2626 818 2734 821
rect 2746 818 2822 821
rect 2826 818 2854 821
rect 2882 818 3838 821
rect 3890 818 4158 821
rect 4170 818 4190 821
rect 4234 818 4286 821
rect 4330 818 4358 821
rect 538 808 582 811
rect 618 808 742 811
rect 874 808 894 811
rect 1066 808 1102 811
rect 1290 808 1406 811
rect 1490 808 1497 811
rect 1642 808 1678 811
rect 1738 808 1806 811
rect 1954 808 2302 811
rect 2610 808 2638 811
rect 2666 808 2678 811
rect 2742 811 2745 818
rect 2690 808 2745 811
rect 2898 808 3318 811
rect 3570 808 4302 811
rect 392 803 394 807
rect 398 803 401 807
rect 406 803 408 807
rect 1416 803 1418 807
rect 1422 803 1425 807
rect 1430 803 1432 807
rect 1494 802 1497 808
rect 1702 802 1705 808
rect 2440 803 2442 807
rect 2446 803 2449 807
rect 2454 803 2456 807
rect 3472 803 3474 807
rect 3478 803 3481 807
rect 3486 803 3488 807
rect 930 798 934 801
rect 1010 798 1310 801
rect 1354 798 1406 801
rect 1642 798 1646 801
rect 1866 798 2078 801
rect 2082 798 2414 801
rect 2466 798 2662 801
rect 2674 798 2678 801
rect 2682 798 2814 801
rect 2890 798 3038 801
rect 3170 798 3206 801
rect 3210 798 3222 801
rect 3498 798 3646 801
rect 3786 798 3894 801
rect 3930 798 4054 801
rect 4066 798 4126 801
rect -26 791 -22 792
rect -26 788 38 791
rect 390 788 534 791
rect 730 788 734 791
rect 1330 788 1422 791
rect 1594 788 3046 791
rect 3050 788 3246 791
rect 3258 788 3294 791
rect 3994 788 4022 791
rect 4026 788 4118 791
rect 390 782 393 788
rect 106 778 230 781
rect 426 778 430 781
rect 434 778 734 781
rect 810 778 934 781
rect 1210 778 1262 781
rect 1614 778 1622 781
rect 1626 778 1862 781
rect 1866 778 2038 781
rect 2162 778 2206 781
rect 2298 778 2302 781
rect 2306 778 2430 781
rect 2506 778 2558 781
rect 2778 778 2878 781
rect 3050 778 3118 781
rect 3122 778 3350 781
rect 3354 778 3510 781
rect 3514 778 3582 781
rect 3610 778 3654 781
rect 3826 778 3854 781
rect 3858 778 3942 781
rect 4142 778 4238 781
rect -26 771 -22 772
rect 6 771 9 778
rect 1598 772 1601 778
rect -26 768 9 771
rect 26 768 318 771
rect 722 768 758 771
rect 1202 768 1470 771
rect 1562 768 1574 771
rect 1602 768 1686 771
rect 2018 768 2094 771
rect 2274 768 2502 771
rect 2506 768 2574 771
rect 2610 768 2638 771
rect 2654 768 2662 771
rect 2666 768 2846 771
rect 2858 768 3134 771
rect 3298 768 3526 771
rect 3618 768 3622 771
rect 3658 768 3662 771
rect 3714 768 3726 771
rect 3730 768 3742 771
rect 3850 768 3870 771
rect 3930 768 3934 771
rect 3962 768 4006 771
rect 4010 768 4030 771
rect 4050 768 4054 771
rect 4142 771 4145 778
rect 4106 768 4145 771
rect 4278 771 4281 778
rect 4234 768 4310 771
rect -26 758 598 761
rect 602 758 630 761
rect 634 758 774 761
rect 1122 758 1126 761
rect 1138 758 1174 761
rect 1218 758 1254 761
rect 1482 758 1494 761
rect 1530 758 1542 761
rect 1546 758 1726 761
rect 1766 761 1769 768
rect 1730 758 1782 761
rect 2014 761 2017 768
rect 3566 762 3569 768
rect 1890 758 2017 761
rect 2034 758 2038 761
rect 2074 758 2078 761
rect 2194 758 2326 761
rect 2386 758 2390 761
rect 2450 758 2478 761
rect 2498 758 2894 761
rect 2922 758 2966 761
rect 3202 758 3270 761
rect 3274 758 3454 761
rect 3466 758 3494 761
rect 3522 758 3558 761
rect 3590 761 3593 768
rect 3590 758 3606 761
rect 3618 758 3686 761
rect 3690 758 3790 761
rect 3826 758 3830 761
rect 3930 758 3934 761
rect 4002 758 4062 761
rect 4338 758 4374 761
rect -26 752 -23 758
rect 2910 752 2913 758
rect 3806 752 3809 758
rect 4110 752 4113 758
rect 4118 752 4121 758
rect 4198 752 4201 758
rect -26 748 -22 752
rect 530 748 702 751
rect 730 748 734 751
rect 754 748 982 751
rect 1118 748 1126 751
rect 1130 748 1190 751
rect 1306 748 1430 751
rect 1458 748 1462 751
rect 1466 748 1630 751
rect 1634 748 1694 751
rect 1730 748 1734 751
rect 1746 748 1798 751
rect 1858 748 1926 751
rect 1930 748 1966 751
rect 1978 748 2014 751
rect 2018 748 2022 751
rect 2026 748 2038 751
rect 2050 748 2254 751
rect 2354 748 2358 751
rect 2402 748 2438 751
rect 2522 748 2526 751
rect 2570 748 2582 751
rect 2586 748 2638 751
rect 2674 748 2678 751
rect 2930 748 2982 751
rect 3154 748 3281 751
rect 3290 748 3310 751
rect 3386 748 3638 751
rect 3642 748 3646 751
rect 3722 748 3750 751
rect 3826 748 3846 751
rect 3850 748 3854 751
rect 3922 748 3926 751
rect 3954 748 3990 751
rect 4226 748 4254 751
rect 4258 748 4270 751
rect 4274 748 4302 751
rect 4370 748 4382 751
rect 4386 748 4390 751
rect 158 742 161 748
rect 1118 742 1121 748
rect 1702 742 1705 748
rect 274 738 286 741
rect 290 738 342 741
rect 346 738 366 741
rect 570 738 574 741
rect 674 738 726 741
rect 738 738 766 741
rect 838 738 918 741
rect 1178 738 1214 741
rect 1318 738 1334 741
rect 1354 738 1366 741
rect 1466 738 1470 741
rect 1490 738 1494 741
rect 1498 738 1638 741
rect 1674 738 1686 741
rect 1722 738 1766 741
rect 1802 738 1806 741
rect 2002 738 2086 741
rect 2226 738 2230 741
rect 2294 741 2297 748
rect 2294 738 2302 741
rect 2354 738 2358 741
rect 2362 738 2390 741
rect 2402 738 2406 741
rect 2518 738 2582 741
rect 2586 738 2598 741
rect 2610 738 2614 741
rect 2618 738 2654 741
rect 2774 741 2777 748
rect 3278 742 3281 748
rect 4062 742 4065 748
rect 2774 738 2838 741
rect 2866 738 2870 741
rect 3018 738 3038 741
rect 3042 738 3222 741
rect 3298 738 3302 741
rect 3506 738 3598 741
rect 3634 738 3638 741
rect 3794 738 3830 741
rect 3858 738 3910 741
rect 4170 738 4246 741
rect 4250 738 4294 741
rect 838 732 841 738
rect 1070 732 1073 738
rect 1318 732 1321 738
rect 142 728 214 731
rect 562 728 646 731
rect 650 728 662 731
rect 666 728 710 731
rect 722 728 726 731
rect 1082 728 1142 731
rect 1146 728 1246 731
rect 1442 728 1462 731
rect 1498 728 1526 731
rect 1614 728 1622 731
rect 1634 728 1838 731
rect 1842 728 1894 731
rect 1922 728 1950 731
rect 1954 728 2014 731
rect 2158 731 2161 738
rect 2082 728 2161 731
rect 2174 732 2177 738
rect 2250 728 2281 731
rect 142 722 145 728
rect 854 722 857 728
rect 1614 722 1617 728
rect 1002 718 1110 721
rect 1154 718 1438 721
rect 1474 718 1518 721
rect 1530 718 1574 721
rect 1658 718 1662 721
rect 1730 718 1806 721
rect 1834 718 1838 721
rect 1894 721 1897 728
rect 2278 722 2281 728
rect 2510 731 2513 738
rect 2506 728 2513 731
rect 2518 732 2521 738
rect 2758 732 2761 738
rect 2530 728 2534 731
rect 2562 728 2654 731
rect 2714 728 2750 731
rect 2914 728 2926 731
rect 2930 728 2998 731
rect 3002 728 3110 731
rect 3422 728 3534 731
rect 3538 728 3542 731
rect 3562 728 3590 731
rect 3618 728 3702 731
rect 3742 731 3745 738
rect 3714 728 3782 731
rect 3802 728 3862 731
rect 3890 728 3910 731
rect 4034 728 4094 731
rect 4098 728 4126 731
rect 4130 728 4342 731
rect 1894 718 1998 721
rect 2010 718 2038 721
rect 2042 718 2158 721
rect 2162 718 2190 721
rect 2286 721 2289 728
rect 2550 722 2553 728
rect 2286 718 2518 721
rect 2722 718 2726 721
rect 2982 718 2990 721
rect 2994 718 3014 721
rect 3074 718 3094 721
rect 3178 718 3302 721
rect 3310 721 3313 728
rect 3422 722 3425 728
rect 3310 718 3422 721
rect 3522 718 4014 721
rect 4194 718 4214 721
rect 1646 712 1649 718
rect 1814 712 1817 718
rect 170 708 222 711
rect 226 708 302 711
rect 442 708 478 711
rect 658 708 678 711
rect 682 708 702 711
rect 706 708 878 711
rect 1242 708 1390 711
rect 1394 708 1422 711
rect 1434 708 1494 711
rect 1506 708 1606 711
rect 1618 708 1638 711
rect 1658 708 1662 711
rect 1874 708 1910 711
rect 2006 711 2009 718
rect 1978 708 2009 711
rect 2114 708 2366 711
rect 2426 708 2470 711
rect 2474 708 2590 711
rect 2602 708 2614 711
rect 2698 708 2726 711
rect 2730 708 2822 711
rect 2826 708 2878 711
rect 2978 708 3134 711
rect 3250 708 3966 711
rect 4162 708 4230 711
rect 896 703 898 707
rect 902 703 905 707
rect 910 703 912 707
rect 1928 703 1930 707
rect 1934 703 1937 707
rect 1942 703 1944 707
rect 2952 703 2954 707
rect 2958 703 2961 707
rect 2966 703 2968 707
rect 3976 703 3978 707
rect 3982 703 3985 707
rect 3990 703 3992 707
rect 314 698 422 701
rect 442 698 454 701
rect 458 698 470 701
rect 474 698 590 701
rect 626 698 710 701
rect 922 698 1038 701
rect 1082 698 1086 701
rect 1106 698 1134 701
rect 1202 698 1238 701
rect 1298 698 1326 701
rect 1402 698 1558 701
rect 1570 698 1654 701
rect 1658 698 1694 701
rect 2090 698 2134 701
rect 2186 698 2190 701
rect 2314 698 2318 701
rect 2490 698 2526 701
rect 2530 698 2606 701
rect 2610 698 2846 701
rect 2994 698 3126 701
rect 3234 698 3334 701
rect 3338 698 3358 701
rect 3418 698 3422 701
rect 3442 698 3694 701
rect 3698 698 3742 701
rect 3770 698 3798 701
rect 3850 698 3870 701
rect 3874 698 3902 701
rect 1846 692 1849 698
rect 234 688 254 691
rect 258 688 534 691
rect 650 688 769 691
rect 522 678 582 681
rect 630 681 633 688
rect 766 682 769 688
rect 958 688 1078 691
rect 1082 688 1094 691
rect 1250 688 1334 691
rect 1450 688 1774 691
rect 1778 688 1782 691
rect 1794 688 1822 691
rect 1906 688 2190 691
rect 2194 688 2286 691
rect 2290 688 2318 691
rect 2330 688 2374 691
rect 2626 688 2630 691
rect 2650 688 2694 691
rect 2698 688 2894 691
rect 2970 688 3022 691
rect 3242 688 3262 691
rect 3270 688 3342 691
rect 3346 688 3358 691
rect 3370 688 3398 691
rect 3410 688 3414 691
rect 3690 688 4014 691
rect 4054 688 4206 691
rect 958 682 961 688
rect 3270 682 3273 688
rect 586 678 633 681
rect 778 678 886 681
rect 1114 678 1374 681
rect 1386 678 1438 681
rect 1458 678 1470 681
rect 1498 678 1566 681
rect 1570 678 1598 681
rect 1706 678 1750 681
rect 1786 678 1822 681
rect 1826 678 1870 681
rect 1882 678 1886 681
rect 1930 678 1982 681
rect 2138 678 2302 681
rect 2306 678 2350 681
rect 2546 678 2622 681
rect 2634 678 2662 681
rect 2674 678 2790 681
rect 2802 678 2854 681
rect 2938 678 2958 681
rect 2966 678 3022 681
rect 3258 678 3270 681
rect 3546 678 3558 681
rect 3590 681 3593 688
rect 3562 678 3593 681
rect 3630 682 3633 688
rect 3682 678 3718 681
rect 3722 678 3750 681
rect 3774 678 3862 681
rect 4054 681 4057 688
rect 3882 678 4057 681
rect 4178 678 4238 681
rect 4242 678 4382 681
rect 134 672 137 678
rect 382 672 385 678
rect 202 668 326 671
rect 470 671 473 678
rect 470 668 510 671
rect 646 671 649 678
rect 646 668 694 671
rect 722 668 750 671
rect 774 671 777 678
rect 1446 672 1449 678
rect 1486 672 1489 678
rect 754 668 777 671
rect 818 668 838 671
rect 1034 668 1126 671
rect 1234 668 1238 671
rect 1242 668 1278 671
rect 1466 668 1478 671
rect 1610 668 1881 671
rect 1898 668 1942 671
rect 1946 668 2046 671
rect 2094 671 2097 678
rect 2094 668 2110 671
rect 2202 668 2230 671
rect 2502 671 2505 678
rect 2402 668 2505 671
rect 2618 668 2758 671
rect 2802 668 2886 671
rect 2914 668 2918 671
rect 2966 671 2969 678
rect 3774 672 3777 678
rect 2922 668 2969 671
rect 2978 668 3006 671
rect 3010 668 3070 671
rect 3306 668 3334 671
rect 3338 668 3374 671
rect 3378 668 3686 671
rect 3706 668 3774 671
rect 3810 668 3838 671
rect 3870 671 3873 678
rect 3842 668 3873 671
rect 3878 672 3881 678
rect 4026 668 4086 671
rect 4130 668 4142 671
rect 4202 668 4310 671
rect 4314 668 4334 671
rect 4362 668 4374 671
rect 194 658 230 661
rect 826 658 846 661
rect 858 658 950 661
rect 974 661 977 668
rect 954 658 977 661
rect 1002 658 1022 661
rect 1042 658 1166 661
rect 1218 658 1265 661
rect 1290 658 1310 661
rect 1430 661 1433 668
rect 1402 658 1433 661
rect 1494 661 1497 668
rect 1518 662 1521 668
rect 1606 662 1609 668
rect 1458 658 1510 661
rect 1618 658 1622 661
rect 1674 658 1678 661
rect 1738 658 1742 661
rect 1762 658 1790 661
rect 1878 661 1881 668
rect 2310 662 2313 668
rect 1878 658 1894 661
rect 1898 658 1958 661
rect 1978 658 2158 661
rect 2226 658 2289 661
rect 2338 658 2350 661
rect 2586 658 2606 661
rect 2610 658 2662 661
rect 2722 658 2750 661
rect 2794 658 2830 661
rect 2950 658 2990 661
rect 3002 658 3006 661
rect 3042 658 3062 661
rect 3362 658 3366 661
rect 3394 658 3398 661
rect 3458 658 3470 661
rect 3486 658 3494 661
rect 3514 658 3550 661
rect 3674 658 3718 661
rect 3722 658 3750 661
rect 3778 658 3782 661
rect 3786 658 3798 661
rect 3866 658 3886 661
rect 4038 658 4046 661
rect 4050 658 4054 661
rect 4102 661 4105 668
rect 4102 658 4118 661
rect 4218 658 4222 661
rect 4282 658 4318 661
rect 4322 658 4350 661
rect -26 651 -22 652
rect -26 648 6 651
rect 714 648 838 651
rect 842 648 926 651
rect 974 651 977 658
rect 1262 652 1265 658
rect 2286 652 2289 658
rect 2950 652 2953 658
rect 974 648 1214 651
rect 1226 648 1230 651
rect 1250 648 1254 651
rect 1314 648 1318 651
rect 1466 648 1478 651
rect 1498 648 1566 651
rect 1590 648 1670 651
rect 1674 648 1718 651
rect 1730 648 1758 651
rect 1882 648 2262 651
rect 2298 648 2342 651
rect 2378 648 2630 651
rect 2762 648 2801 651
rect 2826 648 2838 651
rect 2986 648 2990 651
rect 3006 648 3214 651
rect 3258 648 3262 651
rect 3290 648 3382 651
rect 3406 648 3414 651
rect 3486 651 3489 658
rect 3614 652 3617 658
rect 3418 648 3489 651
rect 3494 648 3526 651
rect 3546 648 3566 651
rect 3754 648 3774 651
rect 3822 651 3825 658
rect 3822 648 3846 651
rect 3898 648 3902 651
rect 4006 651 4009 658
rect 4006 648 4070 651
rect 4178 648 4262 651
rect 4298 648 4302 651
rect 1590 642 1593 648
rect 1766 642 1769 648
rect 2798 642 2801 648
rect 3006 642 3009 648
rect 3494 642 3497 648
rect 4078 642 4081 648
rect 786 638 982 641
rect 1026 638 1030 641
rect 1082 638 1422 641
rect 1490 638 1526 641
rect 1658 638 1686 641
rect 1698 638 1710 641
rect 1714 638 1742 641
rect 2210 638 2214 641
rect 2234 638 2238 641
rect 2258 638 2310 641
rect 2314 638 2350 641
rect 2418 638 2630 641
rect 2634 638 2638 641
rect 3226 638 3417 641
rect 3458 638 3494 641
rect 3506 638 3646 641
rect 3650 638 3830 641
rect 3970 638 3982 641
rect 4010 638 4046 641
rect 4066 638 4070 641
rect 4090 638 4166 641
rect 4298 638 4310 641
rect 4330 638 4342 641
rect 114 628 118 631
rect 138 628 1017 631
rect 1210 628 1270 631
rect 1334 628 1502 631
rect 1522 628 1574 631
rect 2266 628 2902 631
rect 2914 628 2998 631
rect 3082 628 3110 631
rect 3114 628 3350 631
rect 3414 631 3417 638
rect 3414 628 3558 631
rect 3578 628 3809 631
rect 3978 628 4054 631
rect 4066 628 4142 631
rect 1014 622 1017 628
rect 1334 622 1337 628
rect 3806 622 3809 628
rect 122 618 270 621
rect 282 618 286 621
rect 1122 618 1198 621
rect 1202 618 1334 621
rect 1426 618 1638 621
rect 1642 618 1926 621
rect 2354 618 2758 621
rect 2762 618 3598 621
rect 3602 618 3686 621
rect 4138 618 4206 621
rect 4210 618 4262 621
rect 98 608 150 611
rect 938 608 1366 611
rect 1594 608 1646 611
rect 2026 608 2158 611
rect 2242 608 2278 611
rect 2282 608 2422 611
rect 2482 608 2502 611
rect 2658 608 2790 611
rect 2794 608 3230 611
rect 3242 608 3374 611
rect 3410 608 3430 611
rect 3554 608 3598 611
rect 3642 608 3678 611
rect 3714 608 3958 611
rect 4274 608 4366 611
rect 392 603 394 607
rect 398 603 401 607
rect 406 603 408 607
rect 1416 603 1418 607
rect 1422 603 1425 607
rect 1430 603 1432 607
rect 2440 603 2442 607
rect 2446 603 2449 607
rect 2454 603 2456 607
rect 3472 603 3474 607
rect 3478 603 3481 607
rect 3486 603 3488 607
rect 970 598 1118 601
rect 1130 598 1142 601
rect 1442 598 1974 601
rect 2002 598 2166 601
rect 2386 598 2422 601
rect 2490 598 2494 601
rect 2538 598 2750 601
rect 2778 598 3350 601
rect 3570 598 4270 601
rect 626 588 782 591
rect 810 588 838 591
rect 1082 588 1086 591
rect 1310 588 1734 591
rect 1738 588 1910 591
rect 1922 588 1942 591
rect 1978 588 2142 591
rect 2226 588 2318 591
rect 2426 588 2446 591
rect 2450 588 2574 591
rect 2594 588 2854 591
rect 2890 588 2894 591
rect 2898 588 3062 591
rect 3090 588 3158 591
rect 3162 588 3198 591
rect 3218 588 3286 591
rect 3306 588 3334 591
rect 3442 588 3566 591
rect 3602 588 3614 591
rect 3722 588 3726 591
rect 3802 588 3934 591
rect 1310 582 1313 588
rect 282 578 438 581
rect 634 578 998 581
rect 1362 578 1374 581
rect 1442 578 1678 581
rect 1682 578 1910 581
rect 1914 578 2246 581
rect 2410 578 2542 581
rect 2690 578 2734 581
rect 2738 578 2774 581
rect 2778 578 2878 581
rect 3070 581 3073 588
rect 3070 578 3174 581
rect 3178 578 3566 581
rect 3594 578 3654 581
rect 3682 578 3790 581
rect 4034 578 4038 581
rect 4042 578 4062 581
rect 4066 578 4094 581
rect 4102 581 4105 588
rect 4102 578 4246 581
rect 410 568 414 571
rect 802 568 814 571
rect 1382 571 1385 578
rect 986 568 1385 571
rect 1394 568 1406 571
rect 1450 568 1462 571
rect 1506 568 1510 571
rect 1514 568 1534 571
rect 1538 568 1630 571
rect 1634 568 1638 571
rect 1666 568 1694 571
rect 1714 568 1782 571
rect 1802 568 1846 571
rect 1866 568 1921 571
rect 1938 568 1974 571
rect 1994 568 2022 571
rect 2042 568 2102 571
rect 2118 568 2174 571
rect 2186 568 2206 571
rect 2282 568 2350 571
rect 2394 568 2649 571
rect 2658 568 2782 571
rect 2786 568 3254 571
rect 3314 568 3326 571
rect 3330 568 3518 571
rect 3538 568 3574 571
rect 3578 568 3702 571
rect 3810 568 3894 571
rect 3914 568 3942 571
rect 3946 568 3958 571
rect 3962 568 3990 571
rect 3994 568 4086 571
rect 4106 568 4134 571
rect 4138 568 4158 571
rect 4234 568 4278 571
rect 4282 568 4310 571
rect 4346 568 4374 571
rect 1918 562 1921 568
rect 2118 562 2121 568
rect 154 558 438 561
rect 450 558 542 561
rect 546 558 870 561
rect 1090 558 1094 561
rect 1130 558 1270 561
rect 1330 558 1609 561
rect 1618 558 1742 561
rect 1794 558 1806 561
rect 1986 558 2118 561
rect 2154 558 2206 561
rect 2222 561 2225 568
rect 2646 562 2649 568
rect 2210 558 2225 561
rect 2330 558 2398 561
rect 2594 558 2606 561
rect 2610 558 2614 561
rect 2650 558 2670 561
rect 2682 558 2686 561
rect 2714 558 2718 561
rect 2826 558 2830 561
rect 3130 558 3166 561
rect 3170 558 3174 561
rect 3194 558 3230 561
rect 3234 558 3278 561
rect 3338 558 3342 561
rect 3618 558 3718 561
rect 3722 558 3774 561
rect 3806 561 3809 568
rect 4190 562 4193 568
rect 3794 558 3809 561
rect 3882 558 3894 561
rect 3922 558 3950 561
rect 3954 558 3966 561
rect 4074 558 4078 561
rect 4106 558 4110 561
rect 4138 558 4142 561
rect 4178 558 4182 561
rect 4258 558 4326 561
rect 4330 558 4334 561
rect 186 548 190 551
rect 434 548 582 551
rect 850 548 862 551
rect 866 548 958 551
rect 962 548 974 551
rect 1050 548 1110 551
rect 1114 548 1158 551
rect 1282 548 1286 551
rect 1394 548 1406 551
rect 1418 548 1422 551
rect 1458 548 1478 551
rect 1482 548 1502 551
rect 1506 548 1534 551
rect 1570 548 1598 551
rect 1606 551 1609 558
rect 3118 552 3121 558
rect 1606 548 1662 551
rect 1690 548 1774 551
rect 1778 548 1806 551
rect 1810 548 1814 551
rect 1818 548 1870 551
rect 1898 548 1950 551
rect 1954 548 1958 551
rect 1974 548 2022 551
rect 2026 548 2046 551
rect 2162 548 2214 551
rect 2218 548 2382 551
rect 2386 548 2582 551
rect 2594 548 2622 551
rect 2626 548 2726 551
rect 2746 548 2806 551
rect 2810 548 2926 551
rect 3138 548 3150 551
rect 3154 548 3222 551
rect 3258 548 3302 551
rect 3470 551 3473 558
rect 3902 552 3905 558
rect 3466 548 3473 551
rect 3522 548 3646 551
rect 3650 548 3742 551
rect 3938 548 3982 551
rect 4026 548 4030 551
rect 4034 548 4062 551
rect 4066 548 4078 551
rect 4082 548 4110 551
rect 4114 548 4142 551
rect 4166 551 4169 558
rect 4166 548 4174 551
rect 4194 548 4262 551
rect 4274 548 4278 551
rect 4282 548 4318 551
rect 4354 548 4358 551
rect 18 538 78 541
rect 178 538 422 541
rect 426 538 566 541
rect 570 538 590 541
rect 710 538 806 541
rect 842 538 1102 541
rect 1114 538 1230 541
rect 1290 538 1430 541
rect 1434 538 1446 541
rect 1594 538 1646 541
rect 1650 538 1670 541
rect 1714 538 1726 541
rect 1818 538 1854 541
rect 1974 541 1977 548
rect 1882 538 1977 541
rect 1986 538 1990 541
rect 2162 538 2166 541
rect 2170 538 2206 541
rect 2258 538 2294 541
rect 2322 538 2478 541
rect 2602 538 2614 541
rect 2618 540 2662 541
rect 2666 540 2718 541
rect 2618 538 2718 540
rect 2722 538 2782 541
rect 2786 538 2806 541
rect 2990 541 2993 548
rect 3094 541 3097 548
rect 2990 538 3097 541
rect 3122 538 3174 541
rect 3210 538 3214 541
rect 3242 538 3270 541
rect 3314 538 3638 541
rect 3754 538 3774 541
rect 3874 538 3886 541
rect 4290 538 4294 541
rect 710 532 713 538
rect 1478 532 1481 538
rect 1518 532 1521 538
rect 146 528 150 531
rect 154 528 190 531
rect 194 528 297 531
rect 402 528 566 531
rect 570 528 697 531
rect 1130 528 1214 531
rect 1218 528 1238 531
rect 1378 528 1398 531
rect 1554 528 1558 531
rect 1590 528 1606 531
rect 1626 528 1678 531
rect 1754 528 1758 531
rect 1778 528 1782 531
rect 1810 528 1825 531
rect 1858 528 2006 531
rect 2054 531 2057 538
rect 2026 528 2182 531
rect 2186 528 2334 531
rect 2338 528 2622 531
rect 2750 528 2838 531
rect 2974 531 2977 538
rect 2874 528 2977 531
rect 3210 528 3233 531
rect 3258 528 3310 531
rect 3514 528 3558 531
rect 3562 528 3614 531
rect 3650 528 3822 531
rect 3826 528 3846 531
rect 3922 528 4206 531
rect 4218 528 4270 531
rect 4274 528 4342 531
rect 294 522 297 528
rect 694 522 697 528
rect 722 518 758 521
rect 762 518 782 521
rect 786 518 886 521
rect 890 518 982 521
rect 1170 518 1246 521
rect 1258 518 1302 521
rect 1590 521 1593 528
rect 1822 522 1825 528
rect 2750 522 2753 528
rect 3230 522 3233 528
rect 3422 522 3425 528
rect 1394 518 1593 521
rect 1602 518 1614 521
rect 2026 518 2110 521
rect 2138 518 2262 521
rect 2334 518 2342 521
rect 2346 518 2358 521
rect 2634 518 2662 521
rect 2682 518 2702 521
rect 2778 518 2822 521
rect 2826 518 3198 521
rect 3586 518 4046 521
rect 4210 518 4238 521
rect 922 508 974 511
rect 978 508 998 511
rect 1138 508 1510 511
rect 1514 508 1774 511
rect 2018 508 2030 511
rect 2242 508 2654 511
rect 2674 508 2710 511
rect 3018 508 3246 511
rect 3250 508 3294 511
rect 3306 508 3574 511
rect 3578 508 3582 511
rect 3802 508 3814 511
rect 4002 508 4302 511
rect 896 503 898 507
rect 902 503 905 507
rect 910 503 912 507
rect 1928 503 1930 507
rect 1934 503 1937 507
rect 1942 503 1944 507
rect 2952 503 2954 507
rect 2958 503 2961 507
rect 2966 503 2968 507
rect 3976 503 3978 507
rect 3982 503 3985 507
rect 3990 503 3992 507
rect 698 498 750 501
rect 1074 498 1462 501
rect 1554 498 1742 501
rect 1954 498 2086 501
rect 2090 498 2198 501
rect 2426 498 2550 501
rect 2554 498 2558 501
rect 2562 498 2678 501
rect 2690 498 2758 501
rect 2762 498 2934 501
rect 3166 498 3638 501
rect 3642 498 3953 501
rect 4050 498 4054 501
rect 886 491 889 498
rect 3166 492 3169 498
rect 886 488 934 491
rect 938 488 1014 491
rect 1082 488 1118 491
rect 1146 488 1238 491
rect 1586 488 1638 491
rect 1706 488 1750 491
rect 1758 488 1766 491
rect 1770 488 1830 491
rect 1834 488 1998 491
rect 2042 488 2094 491
rect 2258 488 2262 491
rect 2354 488 2478 491
rect 2482 488 2518 491
rect 2706 488 2798 491
rect 2954 488 2958 491
rect 3062 488 3166 491
rect 3354 488 3406 491
rect 3426 488 3558 491
rect 3650 488 3694 491
rect 3794 488 3814 491
rect 3950 491 3953 498
rect 3950 488 4014 491
rect 4242 488 4270 491
rect 66 478 142 481
rect 286 481 289 488
rect 146 478 289 481
rect 654 481 657 488
rect 862 481 865 488
rect 538 478 865 481
rect 1046 481 1049 488
rect 1270 482 1273 488
rect 2006 482 2009 488
rect 3062 482 3065 488
rect 994 478 1134 481
rect 1218 478 1222 481
rect 1258 478 1262 481
rect 1306 478 1414 481
rect 1458 478 1478 481
rect 1482 478 1486 481
rect 1514 478 1534 481
rect 1538 478 1590 481
rect 1658 478 1710 481
rect 1714 478 1790 481
rect 2058 478 2150 481
rect 2154 478 2158 481
rect 2274 478 2390 481
rect 2550 478 2798 481
rect 2882 478 3062 481
rect 3074 478 3094 481
rect 3114 478 3158 481
rect 3162 478 3166 481
rect 3178 478 3206 481
rect 3406 481 3409 488
rect 3406 478 3550 481
rect 3602 478 3702 481
rect 3770 478 3838 481
rect 3842 478 3854 481
rect 3858 478 3870 481
rect 3874 478 3910 481
rect 3946 478 4006 481
rect 4066 478 4153 481
rect 4162 478 4182 481
rect 4210 478 4294 481
rect 1606 472 1609 478
rect 722 468 742 471
rect 986 468 1110 471
rect 1146 468 1150 471
rect 1186 468 1358 471
rect 1362 468 1446 471
rect 1482 468 1494 471
rect 1570 468 1574 471
rect 1742 468 1814 471
rect 1822 471 1825 478
rect 2550 472 2553 478
rect 1822 468 1838 471
rect 1842 468 1950 471
rect 2002 468 2086 471
rect 2178 468 2374 471
rect 2378 468 2406 471
rect 2514 468 2534 471
rect 2738 468 2766 471
rect 2938 468 2974 471
rect 3042 468 3113 471
rect 3122 468 3126 471
rect 3218 468 3230 471
rect 3306 468 3310 471
rect 3594 468 3598 471
rect 3702 471 3705 478
rect 3702 468 3742 471
rect 3770 468 3782 471
rect 3786 468 3878 471
rect 3898 468 3937 471
rect 4002 468 4006 471
rect 4150 471 4153 478
rect 4150 468 4174 471
rect 4290 468 4310 471
rect 182 461 185 468
rect 1454 462 1457 468
rect 1526 462 1529 468
rect 182 458 230 461
rect 274 458 681 461
rect 714 458 734 461
rect 986 458 1166 461
rect 1370 458 1382 461
rect 1466 458 1478 461
rect 1482 458 1518 461
rect 1582 461 1585 468
rect 1742 462 1745 468
rect 2462 462 2465 468
rect 1582 458 1614 461
rect 1770 458 1782 461
rect 1790 458 1862 461
rect 1866 458 1873 461
rect 1898 458 2342 461
rect 2354 458 2358 461
rect 2490 458 2529 461
rect 2646 461 2649 468
rect 2586 458 2649 461
rect 2770 458 2774 461
rect 3050 458 3054 461
rect 3082 458 3094 461
rect 3110 461 3113 468
rect 3166 462 3169 468
rect 3182 462 3185 468
rect 3110 458 3142 461
rect 3234 458 3238 461
rect 3282 458 3518 461
rect 3602 458 3630 461
rect 3694 461 3697 468
rect 3934 462 3937 468
rect 3674 458 3697 461
rect 3730 458 3774 461
rect 3818 458 3822 461
rect 4038 461 4041 468
rect 4038 458 4054 461
rect 4090 458 4094 461
rect 4102 461 4105 468
rect 4102 458 4150 461
rect 4186 458 4190 461
rect 4246 461 4249 468
rect 4226 458 4249 461
rect 4258 458 4278 461
rect 4346 458 4366 461
rect -26 451 -22 452
rect -26 448 6 451
rect 678 451 681 458
rect 1534 452 1537 458
rect 678 448 993 451
rect 1026 448 1113 451
rect 1130 448 1134 451
rect 1314 448 1334 451
rect 1570 448 1654 451
rect 1734 448 1774 451
rect 1790 451 1793 458
rect 2526 452 2529 458
rect 1790 448 1798 451
rect 1834 448 1838 451
rect 1866 448 1894 451
rect 2034 448 2078 451
rect 2114 448 2118 451
rect 2146 448 2310 451
rect 2330 448 2390 451
rect 2506 448 2510 451
rect 2538 448 2558 451
rect 2562 448 2566 451
rect 2570 448 2577 451
rect 2594 448 2606 451
rect 2930 448 3022 451
rect 3026 448 3030 451
rect 3158 451 3161 458
rect 3158 448 3190 451
rect 3202 448 3598 451
rect 3610 448 3662 451
rect 3826 448 3838 451
rect 3994 448 4054 451
rect 4082 448 4086 451
rect 4122 448 4126 451
rect 4178 448 4310 451
rect 4314 448 4326 451
rect 4338 448 4342 451
rect 990 442 993 448
rect 410 438 414 441
rect 562 438 566 441
rect 674 438 790 441
rect 1058 438 1102 441
rect 1110 441 1113 448
rect 1142 441 1145 448
rect 1734 442 1737 448
rect 1110 438 1145 441
rect 1394 438 1550 441
rect 2126 441 2129 448
rect 3094 442 3097 448
rect 2010 438 2129 441
rect 2154 438 2334 441
rect 2346 438 2518 441
rect 2522 438 2614 441
rect 2690 438 2806 441
rect 3570 438 3646 441
rect 3682 438 3950 441
rect 4034 438 4110 441
rect 4130 438 4142 441
rect 4234 438 4238 441
rect 4242 438 4326 441
rect 4330 438 4374 441
rect 378 428 558 431
rect 1054 431 1057 438
rect 562 428 1057 431
rect 1122 428 1582 431
rect 1646 431 1649 438
rect 4214 432 4217 438
rect 1646 428 2246 431
rect 2370 428 3926 431
rect 3970 428 4094 431
rect 4098 428 4102 431
rect 4106 428 4150 431
rect 4298 428 4302 431
rect 4322 428 4345 431
rect 4342 422 4345 428
rect 122 418 678 421
rect 682 418 798 421
rect 802 418 854 421
rect 882 418 929 421
rect 1018 418 1174 421
rect 1362 418 1366 421
rect 1650 418 2070 421
rect 2086 418 2094 421
rect 2098 418 2102 421
rect 2114 418 2134 421
rect 2138 418 2486 421
rect 3050 418 3254 421
rect 3730 418 3774 421
rect 3842 418 4206 421
rect 90 408 118 411
rect 490 408 918 411
rect 926 411 929 418
rect 926 408 1062 411
rect 1226 408 1230 411
rect 1298 408 1382 411
rect 1610 408 1854 411
rect 1858 408 1878 411
rect 2106 408 2422 411
rect 2466 408 2566 411
rect 2642 408 2726 411
rect 3114 408 3214 411
rect 3498 408 3798 411
rect 392 403 394 407
rect 398 403 401 407
rect 406 403 408 407
rect 1416 403 1418 407
rect 1422 403 1425 407
rect 1430 403 1432 407
rect 2440 403 2442 407
rect 2446 403 2449 407
rect 2454 403 2456 407
rect 3472 403 3474 407
rect 3478 403 3481 407
rect 3486 403 3488 407
rect 578 398 614 401
rect 618 398 766 401
rect 826 398 846 401
rect 954 398 1030 401
rect 1034 398 1094 401
rect 1490 398 1646 401
rect 1674 398 1702 401
rect 1842 398 2238 401
rect 2290 398 2342 401
rect 2586 398 2654 401
rect 2810 398 3214 401
rect 3538 398 3654 401
rect 3746 398 3854 401
rect 3858 398 3894 401
rect 4074 398 4174 401
rect 4178 398 4262 401
rect 782 392 785 398
rect 98 388 214 391
rect 482 388 526 391
rect 538 388 550 391
rect 554 388 686 391
rect 794 388 1134 391
rect 1838 391 1841 398
rect 2766 392 2769 398
rect 4262 392 4265 398
rect 1234 388 1841 391
rect 2026 388 2030 391
rect 2130 388 2134 391
rect 2238 388 2246 391
rect 2250 388 2486 391
rect 2530 388 2638 391
rect 2642 388 2646 391
rect 2650 388 2702 391
rect 3066 388 3086 391
rect 3194 388 3278 391
rect 3330 388 3430 391
rect 3434 388 3678 391
rect 3710 382 3713 388
rect 114 378 814 381
rect 986 378 998 381
rect 1002 378 1326 381
rect 1402 378 1574 381
rect 1578 378 1710 381
rect 1714 378 1798 381
rect 1810 378 1838 381
rect 1842 378 1918 381
rect 1922 378 1998 381
rect 2106 378 2462 381
rect 2466 378 2558 381
rect 2562 378 2654 381
rect 2658 378 2830 381
rect 3082 378 3102 381
rect 3106 378 3174 381
rect 3178 378 3334 381
rect 3338 378 3414 381
rect 3418 378 3630 381
rect 3634 378 3646 381
rect 3674 378 3686 381
rect 3890 378 4270 381
rect 894 371 897 378
rect 394 368 897 371
rect 1146 368 1190 371
rect 1314 368 1318 371
rect 1354 368 1358 371
rect 1362 368 1374 371
rect 1458 368 1494 371
rect 1514 368 1566 371
rect 1698 368 1894 371
rect 2306 368 2334 371
rect 2338 368 2406 371
rect 2410 368 2478 371
rect 2490 368 2510 371
rect 2514 368 2521 371
rect 2530 368 2534 371
rect 2574 368 2718 371
rect 2722 368 3798 371
rect 3806 368 3814 371
rect 3818 368 3838 371
rect 3854 368 3857 378
rect 4358 372 4361 378
rect 3866 368 3878 371
rect 3938 368 3942 371
rect 4202 368 4230 371
rect 4234 368 4262 371
rect 4266 368 4294 371
rect 4298 368 4326 371
rect 4330 368 4358 371
rect 186 358 302 361
rect 306 358 646 361
rect 974 361 977 368
rect 946 358 977 361
rect 1038 358 1046 361
rect 1050 358 1070 361
rect 1074 358 1094 361
rect 1238 361 1241 368
rect 1194 358 1241 361
rect 1286 361 1289 368
rect 2006 362 2009 368
rect 2574 362 2577 368
rect 1286 358 1318 361
rect 1338 358 1422 361
rect 1474 358 1510 361
rect 1530 358 1542 361
rect 1594 358 1854 361
rect 1986 358 2006 361
rect 2058 358 2230 361
rect 2234 358 2254 361
rect 2258 358 2278 361
rect 2314 358 2342 361
rect 2450 358 2574 361
rect 2626 358 2686 361
rect 2898 358 2974 361
rect 2978 358 2990 361
rect 2998 358 3006 361
rect 3010 358 3062 361
rect 3234 358 3270 361
rect 3378 358 3494 361
rect 3642 358 3694 361
rect 3722 358 3846 361
rect 3850 358 4014 361
rect 4066 358 4166 361
rect 4202 358 4206 361
rect 4234 358 4238 361
rect 4290 358 4294 361
rect -26 351 -22 352
rect -26 348 6 351
rect 26 348 102 351
rect 266 348 278 351
rect 282 348 326 351
rect 330 348 334 351
rect 386 348 526 351
rect 530 348 582 351
rect 602 348 614 351
rect 678 351 681 358
rect 1182 352 1185 358
rect 678 348 710 351
rect 906 348 966 351
rect 978 348 1030 351
rect 1034 348 1150 351
rect 1262 351 1265 358
rect 4278 352 4281 358
rect 1202 348 1265 351
rect 1282 348 1558 351
rect 1570 348 1846 351
rect 1898 348 2166 351
rect 2170 348 2262 351
rect 2282 348 2289 351
rect 2298 348 2318 351
rect 2322 348 2390 351
rect 2482 348 2502 351
rect 2522 348 2542 351
rect 2570 348 2574 351
rect 2634 348 2662 351
rect 2706 348 2734 351
rect 3002 348 3054 351
rect 3266 348 3286 351
rect 3330 348 3366 351
rect 3386 348 3390 351
rect 3466 348 3470 351
rect 3610 348 3614 351
rect 3670 348 3822 351
rect 3842 348 3926 351
rect 3930 348 3982 351
rect 4034 348 4102 351
rect 4194 348 4222 351
rect 4226 348 4254 351
rect 4258 348 4278 351
rect 4282 348 4302 351
rect 4306 348 4350 351
rect 18 338 38 341
rect 538 338 590 341
rect 814 341 817 348
rect 886 342 889 348
rect 814 338 865 341
rect 930 338 1054 341
rect 1066 338 1070 341
rect 1130 338 1230 341
rect 1242 338 1350 341
rect 1386 338 1470 341
rect 1498 338 1526 341
rect 1546 338 1550 341
rect 1594 338 1726 341
rect 1734 338 1750 341
rect 1754 338 1886 341
rect 1938 338 1942 341
rect 1946 338 1990 341
rect 1994 338 2046 341
rect 2242 338 2246 341
rect 2250 338 2334 341
rect 2338 338 2366 341
rect 2386 338 2414 341
rect 2598 341 2601 348
rect 2434 338 2601 341
rect 2866 338 2958 341
rect 2974 341 2977 348
rect 2974 338 3014 341
rect 3050 338 3078 341
rect 3250 338 3254 341
rect 3270 338 3278 341
rect 3282 338 3294 341
rect 3298 338 3342 341
rect 3670 341 3673 348
rect 3346 338 3673 341
rect 3682 338 3718 341
rect 3730 338 3734 341
rect 3746 338 3750 341
rect 3826 338 3854 341
rect 3874 338 3894 341
rect 3906 338 3910 341
rect 3962 338 3998 341
rect 206 332 209 338
rect 694 331 697 338
rect 694 328 854 331
rect 862 331 865 338
rect 1086 331 1089 338
rect 862 328 1089 331
rect 1154 328 1206 331
rect 1218 328 1286 331
rect 1298 328 1310 331
rect 1522 328 1542 331
rect 1558 328 1694 331
rect 1734 331 1737 338
rect 1714 328 1737 331
rect 2002 328 2038 331
rect 2042 328 2070 331
rect 2110 331 2113 338
rect 2090 328 2113 331
rect 2122 328 2310 331
rect 2362 328 2374 331
rect 2606 331 2609 338
rect 2498 328 2609 331
rect 2638 331 2641 338
rect 2618 328 2641 331
rect 2702 331 2705 338
rect 2682 328 2705 331
rect 3650 328 3726 331
rect 3886 328 3926 331
rect 3930 328 3934 331
rect 3938 328 3966 331
rect 4086 331 4089 338
rect 3978 328 4350 331
rect 122 318 142 321
rect 502 321 505 328
rect 362 318 505 321
rect 722 318 726 321
rect 850 318 982 321
rect 1090 318 1214 321
rect 1242 318 1246 321
rect 1338 318 1462 321
rect 1558 321 1561 328
rect 1490 318 1561 321
rect 1570 318 1782 321
rect 1810 318 1830 321
rect 1842 318 2262 321
rect 2390 321 2393 328
rect 3518 322 3521 328
rect 2282 318 2393 321
rect 2402 318 2798 321
rect 3242 318 3302 321
rect 3322 318 3390 321
rect 3610 318 3678 321
rect 3690 318 3702 321
rect 3706 318 3774 321
rect 3790 321 3793 328
rect 3886 322 3889 328
rect 3790 318 3886 321
rect 3918 318 4366 321
rect 718 311 721 318
rect 362 308 721 311
rect 922 308 1494 311
rect 1602 308 1758 311
rect 1826 308 1846 311
rect 2130 308 2486 311
rect 2530 308 2678 311
rect 2802 308 2942 311
rect 3338 308 3486 311
rect 3490 308 3590 311
rect 3918 311 3921 318
rect 3594 308 3921 311
rect 3962 308 3966 311
rect 4074 308 4334 311
rect 4370 308 4374 311
rect 782 302 785 308
rect 896 303 898 307
rect 902 303 905 307
rect 910 303 912 307
rect 1928 303 1930 307
rect 1934 303 1937 307
rect 1942 303 1944 307
rect 2952 303 2954 307
rect 2958 303 2961 307
rect 2966 303 2968 307
rect 3976 303 3978 307
rect 3982 303 3985 307
rect 3990 303 3992 307
rect 194 298 406 301
rect 586 298 630 301
rect 634 298 662 301
rect 666 298 758 301
rect 1010 298 1014 301
rect 1098 298 1198 301
rect 1266 298 1270 301
rect 1338 298 1470 301
rect 1474 298 1670 301
rect 1682 298 1814 301
rect 2082 298 2118 301
rect 2162 298 2206 301
rect 2282 298 2382 301
rect 2402 298 2534 301
rect 2538 298 2622 301
rect 2818 298 2838 301
rect 2850 298 2926 301
rect 2930 298 2934 301
rect 3026 298 3054 301
rect 3058 298 3078 301
rect 3082 298 3118 301
rect 3122 298 3310 301
rect 3314 298 3350 301
rect 3354 298 3382 301
rect 3390 298 3502 301
rect 3562 298 3582 301
rect 3738 298 3814 301
rect 3922 298 3966 301
rect 378 288 382 291
rect 538 288 542 291
rect 778 288 838 291
rect 842 288 950 291
rect 1562 288 1670 291
rect 1730 288 1838 291
rect 1930 288 1990 291
rect 2018 288 2086 291
rect 2170 288 2222 291
rect 2266 288 2358 291
rect 2362 288 2366 291
rect 2386 288 2406 291
rect 2570 288 2598 291
rect 2746 288 2806 291
rect 2818 288 2942 291
rect 2962 288 3030 291
rect 3058 288 3070 291
rect 3138 288 3150 291
rect 3390 291 3393 298
rect 3258 288 3393 291
rect 3442 288 3454 291
rect 3494 288 3526 291
rect 3586 288 3609 291
rect 3630 288 3638 291
rect 3642 288 3662 291
rect 3666 288 3742 291
rect 3770 288 3790 291
rect 3794 288 3801 291
rect 3810 288 3982 291
rect 4258 288 4270 291
rect 262 281 265 288
rect 98 278 265 281
rect 518 282 521 288
rect 810 278 854 281
rect 1046 278 1110 281
rect 1122 278 1134 281
rect 1322 278 1518 281
rect 1538 278 1590 281
rect 1610 278 1614 281
rect 1626 278 1638 281
rect 1786 278 1798 281
rect 1866 278 1878 281
rect 2094 281 2097 288
rect 2558 282 2561 288
rect 1882 278 2041 281
rect 2094 278 2126 281
rect 2130 278 2270 281
rect 2450 278 2494 281
rect 2686 281 2689 288
rect 2686 278 2702 281
rect 2942 281 2945 288
rect 3406 282 3409 288
rect 2942 278 3102 281
rect 3146 278 3174 281
rect 3306 278 3334 281
rect 3338 278 3398 281
rect 3414 281 3417 288
rect 3494 282 3497 288
rect 3606 282 3609 288
rect 3414 278 3494 281
rect 3522 278 3574 281
rect 3594 278 3598 281
rect 3626 278 3646 281
rect 3658 278 3694 281
rect 3698 278 3718 281
rect 3722 278 3806 281
rect 3922 278 3926 281
rect 3938 278 4102 281
rect 4198 281 4201 288
rect 4198 278 4262 281
rect 4266 278 4286 281
rect 534 272 537 278
rect 394 268 454 271
rect 458 268 478 271
rect 634 268 638 271
rect 670 271 673 278
rect 1046 272 1049 278
rect 670 268 814 271
rect 818 268 825 271
rect 834 268 918 271
rect 1174 271 1177 278
rect 1230 272 1233 278
rect 2038 272 2041 278
rect 1066 268 1177 271
rect 1186 268 1214 271
rect 1234 268 1278 271
rect 1298 268 1374 271
rect 1378 268 1382 271
rect 1402 268 1438 271
rect 1442 268 1446 271
rect 1506 268 1518 271
rect 1530 268 1574 271
rect 1578 268 1814 271
rect 1834 268 1982 271
rect 1994 268 2022 271
rect 2042 268 2070 271
rect 2074 268 2134 271
rect 2138 268 2142 271
rect 2146 268 2206 271
rect 2210 268 2262 271
rect 2310 271 2313 278
rect 2806 272 2809 278
rect 2266 268 2313 271
rect 2370 268 2374 271
rect 2482 268 2518 271
rect 2546 268 2590 271
rect 2738 268 2790 271
rect 2938 268 3062 271
rect 3066 268 3110 271
rect 3162 268 3318 271
rect 3402 268 3566 271
rect 3570 268 3806 271
rect 3810 268 3894 271
rect 3898 268 3926 271
rect 3930 268 4006 271
rect 4082 268 4086 271
rect 4182 271 4185 278
rect 4178 268 4185 271
rect 110 262 113 268
rect 154 258 190 261
rect 418 258 422 261
rect 830 261 833 268
rect 826 258 833 261
rect 906 258 950 261
rect 1034 258 1118 261
rect 1210 258 1246 261
rect 1294 258 1302 261
rect 1306 258 1350 261
rect 1386 258 1406 261
rect 1434 258 1462 261
rect 1486 261 1489 268
rect 1474 258 1489 261
rect 1498 258 1502 261
rect 1506 258 1550 261
rect 1554 258 1790 261
rect 1794 258 1870 261
rect 2034 258 2398 261
rect 2474 258 2510 261
rect 2754 258 2774 261
rect 3058 258 3078 261
rect 3094 258 3134 261
rect 3178 258 3342 261
rect 3378 258 3542 261
rect 3562 258 3590 261
rect 3594 258 3614 261
rect 3682 258 3726 261
rect 3762 258 3793 261
rect 3802 258 3870 261
rect 3890 258 3894 261
rect 3914 258 3934 261
rect 4002 258 4014 261
rect 4050 258 4081 261
rect 4226 258 4286 261
rect 4306 258 4334 261
rect 690 248 838 251
rect 1198 251 1201 258
rect 3094 252 3097 258
rect 3790 252 3793 258
rect 4078 252 4081 258
rect 970 248 1201 251
rect 1218 248 1230 251
rect 1286 248 1294 251
rect 1298 248 1310 251
rect 1354 248 1478 251
rect 1482 248 1526 251
rect 1594 248 1598 251
rect 1722 248 2150 251
rect 2154 248 2230 251
rect 2282 248 2286 251
rect 2330 248 2334 251
rect 2354 248 2358 251
rect 2410 248 2414 251
rect 2430 248 2438 251
rect 2442 248 2478 251
rect 2514 248 2702 251
rect 2866 248 2870 251
rect 3106 248 3134 251
rect 3138 248 3238 251
rect 3370 248 3470 251
rect 3482 248 3502 251
rect 3570 248 3598 251
rect 3634 248 3638 251
rect 3714 248 3742 251
rect 3794 248 3950 251
rect 3954 248 4014 251
rect 862 241 865 248
rect 250 238 865 241
rect 1170 238 1326 241
rect 1330 238 1614 241
rect 2350 241 2353 248
rect 1618 238 2353 241
rect 2410 238 2510 241
rect 2514 238 2822 241
rect 2826 238 3046 241
rect 3050 238 3054 241
rect 3066 238 3846 241
rect 3850 238 3918 241
rect 3986 238 4038 241
rect 362 228 614 231
rect 834 228 894 231
rect 1162 228 1230 231
rect 1234 228 1262 231
rect 1266 228 1350 231
rect 1354 228 1358 231
rect 1362 228 1438 231
rect 1442 228 1454 231
rect 1474 228 1478 231
rect 1554 228 1662 231
rect 1786 228 1886 231
rect 1946 228 2046 231
rect 2098 228 2118 231
rect 2122 228 2182 231
rect 2242 228 2462 231
rect 2466 228 2550 231
rect 2554 228 2590 231
rect 2594 228 3142 231
rect 3242 228 3726 231
rect 3730 228 3766 231
rect 3826 228 3830 231
rect 3898 228 3902 231
rect 4002 228 4070 231
rect 4074 228 4110 231
rect 4114 228 4118 231
rect 4266 228 4294 231
rect 354 218 614 221
rect 858 218 1030 221
rect 1034 218 1110 221
rect 1122 218 1310 221
rect 1386 218 1390 221
rect 1426 218 1486 221
rect 1530 218 1566 221
rect 1662 221 1665 228
rect 1662 218 1838 221
rect 1842 218 2014 221
rect 2042 218 2086 221
rect 2090 218 2134 221
rect 2138 218 2462 221
rect 2466 218 2502 221
rect 2530 218 2854 221
rect 2858 218 3110 221
rect 3114 218 3518 221
rect 3522 218 3542 221
rect 3642 218 3702 221
rect 3706 218 3710 221
rect 3870 221 3873 228
rect 3722 218 3873 221
rect 3890 218 4030 221
rect 678 212 681 218
rect 418 208 438 211
rect 882 208 894 211
rect 906 208 950 211
rect 954 208 1094 211
rect 1206 208 1366 211
rect 1442 208 1646 211
rect 1898 208 2054 211
rect 2058 208 2118 211
rect 2754 208 2830 211
rect 2946 208 2950 211
rect 2978 208 2990 211
rect 3562 208 3710 211
rect 3722 208 3726 211
rect 3738 208 3750 211
rect 3834 208 4046 211
rect 4202 208 4214 211
rect 392 203 394 207
rect 398 203 401 207
rect 406 203 408 207
rect 794 198 1062 201
rect 1206 201 1209 208
rect 1416 203 1418 207
rect 1422 203 1425 207
rect 1430 203 1432 207
rect 2440 203 2442 207
rect 2446 203 2449 207
rect 2454 203 2456 207
rect 2462 202 2465 208
rect 3472 203 3474 207
rect 3478 203 3481 207
rect 3486 203 3488 207
rect 1066 198 1209 201
rect 1218 198 1398 201
rect 1450 198 1582 201
rect 1746 198 2174 201
rect 2290 198 2302 201
rect 2498 198 2542 201
rect 2586 198 2646 201
rect 2722 198 2838 201
rect 2842 198 3358 201
rect 3682 198 3894 201
rect 3906 198 4086 201
rect 2262 192 2265 198
rect 42 188 54 191
rect 58 188 78 191
rect 322 188 790 191
rect 938 188 1078 191
rect 1090 188 1166 191
rect 1194 188 1198 191
rect 1218 188 1249 191
rect 1258 188 1302 191
rect 1322 188 1398 191
rect 1402 188 1462 191
rect 1466 188 2230 191
rect 2426 188 2998 191
rect 3218 188 3246 191
rect 3458 188 3630 191
rect 3658 188 3774 191
rect 3806 188 3918 191
rect 1246 182 1249 188
rect 314 178 374 181
rect 946 178 1238 181
rect 1266 178 1334 181
rect 1498 178 1590 181
rect 1634 178 2006 181
rect 2014 178 2022 181
rect 2026 178 2198 181
rect 2202 178 2326 181
rect 2402 178 2470 181
rect 2474 178 2502 181
rect 2530 178 2534 181
rect 2570 178 2590 181
rect 2610 178 2630 181
rect 2658 178 2662 181
rect 2666 178 2726 181
rect 2730 178 3118 181
rect 3202 178 3406 181
rect 3806 181 3809 188
rect 3410 178 3809 181
rect 3818 178 3862 181
rect 3898 178 3966 181
rect 4274 178 4294 181
rect 4338 178 4342 181
rect 830 171 833 178
rect 738 168 833 171
rect 850 168 966 171
rect 978 168 1014 171
rect 1058 168 1086 171
rect 1114 168 1190 171
rect 1242 168 2254 171
rect 2258 168 2718 171
rect 2874 168 3422 171
rect 3466 168 3470 171
rect 3474 168 3622 171
rect 3670 168 4062 171
rect 4074 168 4110 171
rect 4206 171 4209 178
rect 4114 168 4209 171
rect 4290 168 4390 171
rect 346 158 358 161
rect 810 158 822 161
rect 898 158 934 161
rect 946 158 982 161
rect 1038 161 1041 168
rect 3670 162 3673 168
rect 994 158 1041 161
rect 1082 158 1134 161
rect 1138 158 1182 161
rect 1186 158 1230 161
rect 1250 158 1262 161
rect 1266 158 1270 161
rect 1306 158 1326 161
rect 1338 158 1390 161
rect 1458 158 1494 161
rect 1522 158 1534 161
rect 1570 158 1590 161
rect 1930 158 1934 161
rect 1954 158 2038 161
rect 2058 158 2126 161
rect 2130 158 2190 161
rect 2362 158 2686 161
rect 2690 158 3062 161
rect 3362 158 3670 161
rect 3842 158 3854 161
rect 3882 158 3905 161
rect 3918 158 3926 161
rect 3930 158 3934 161
rect 4042 158 4262 161
rect 4306 158 4318 161
rect 4330 158 4358 161
rect 4362 158 4366 161
rect 218 148 222 151
rect 586 148 630 151
rect 830 148 846 151
rect 906 148 974 151
rect 986 148 1014 151
rect 1018 148 1374 151
rect 1402 148 1406 151
rect 1418 148 1465 151
rect 1530 148 1550 151
rect 1598 151 1601 158
rect 1562 148 1601 151
rect 1618 148 1622 151
rect 1906 148 1958 151
rect 1962 148 2038 151
rect 2050 148 2062 151
rect 2066 148 2073 151
rect 2082 148 2110 151
rect 2146 148 2174 151
rect 2186 148 2286 151
rect 2290 148 2558 151
rect 2562 148 2694 151
rect 2706 148 2710 151
rect 2722 148 3126 151
rect 3394 148 3414 151
rect 3734 151 3737 158
rect 3618 148 3737 151
rect 3814 152 3817 158
rect 3902 152 3905 158
rect 3818 148 3846 151
rect 3978 148 4006 151
rect 4010 148 4142 151
rect 4298 148 4302 151
rect -26 141 -22 142
rect 6 141 9 148
rect 494 142 497 148
rect 694 142 697 148
rect 830 142 833 148
rect -26 138 254 141
rect 834 138 958 141
rect 994 138 1017 141
rect 1026 138 1030 141
rect 1042 138 1110 141
rect 1130 138 1142 141
rect 1154 138 1158 141
rect 1202 138 1246 141
rect 1258 138 1310 141
rect 1378 138 1454 141
rect 1462 141 1465 148
rect 2118 142 2121 148
rect 1462 138 1534 141
rect 1586 138 1614 141
rect 1642 138 1646 141
rect 1650 138 1718 141
rect 1834 138 1894 141
rect 2026 138 2062 141
rect 2066 138 2070 141
rect 2082 138 2086 141
rect 2178 138 2214 141
rect 2218 138 2222 141
rect 2234 138 2414 141
rect 2434 138 2438 141
rect 2466 138 2494 141
rect 2506 138 2646 141
rect 2650 138 2742 141
rect 2746 138 2774 141
rect 2914 138 2934 141
rect 2938 138 2958 141
rect 3058 138 3182 141
rect 3186 138 3286 141
rect 3302 141 3305 148
rect 3926 142 3929 148
rect 3302 138 3358 141
rect 3378 138 3422 141
rect 3618 138 3838 141
rect 3866 138 3878 141
rect 3882 138 3918 141
rect 3950 138 4129 141
rect 4194 138 4318 141
rect 146 128 233 131
rect 866 128 998 131
rect 1014 131 1017 138
rect 1070 132 1073 138
rect 1318 132 1321 138
rect 1726 132 1729 138
rect 1014 128 1038 131
rect 1090 128 1094 131
rect 1122 128 1134 131
rect 1138 128 1286 131
rect 1370 128 1406 131
rect 1418 128 1438 131
rect 1570 128 1710 131
rect 1802 128 1974 131
rect 1998 131 2001 138
rect 3950 132 3953 138
rect 4126 132 4129 138
rect 1998 128 2014 131
rect 2050 128 2350 131
rect 2362 128 2486 131
rect 2546 128 2550 131
rect 2562 128 2566 131
rect 2578 128 2614 131
rect 2642 128 2681 131
rect 2770 128 2854 131
rect 3146 128 3246 131
rect 3442 128 3654 131
rect 3738 128 3742 131
rect 3802 128 3942 131
rect 4314 128 4318 131
rect 4322 128 4374 131
rect 230 122 233 128
rect 618 118 878 121
rect 882 118 1334 121
rect 1346 118 1382 121
rect 1626 118 1654 121
rect 1658 118 1814 121
rect 1974 121 1977 128
rect 2342 122 2345 128
rect 2678 122 2681 128
rect 4302 122 4305 128
rect 1974 118 2006 121
rect 2050 118 2094 121
rect 2098 118 2214 121
rect 2538 118 2590 121
rect 2874 118 3174 121
rect 3186 118 3558 121
rect 3562 118 3662 121
rect 3722 118 3790 121
rect 3810 118 3838 121
rect 4106 118 4262 121
rect 234 108 286 111
rect 642 108 814 111
rect 818 108 870 111
rect 1042 108 1286 111
rect 1330 108 1406 111
rect 1602 108 1806 111
rect 2322 108 2334 111
rect 2354 108 2358 111
rect 2546 108 2638 111
rect 3178 108 3430 111
rect 3434 108 3809 111
rect 4042 108 4086 111
rect 4098 108 4134 111
rect 4138 108 4174 111
rect 4178 108 4350 111
rect 896 103 898 107
rect 902 103 905 107
rect 910 103 912 107
rect 1928 103 1930 107
rect 1934 103 1937 107
rect 1942 103 1944 107
rect 170 98 198 101
rect 570 98 574 101
rect 770 98 774 101
rect 942 98 1358 101
rect 1386 98 1478 101
rect 1522 98 1622 101
rect 1706 98 1726 101
rect 1738 98 1918 101
rect 2010 98 2158 101
rect 2334 101 2337 108
rect 2952 103 2954 107
rect 2958 103 2961 107
rect 2966 103 2968 107
rect 3806 102 3809 108
rect 3976 103 3978 107
rect 3982 103 3985 107
rect 3990 103 3992 107
rect 2334 98 2702 101
rect 2794 98 2806 101
rect 3070 98 3366 101
rect 3378 98 3454 101
rect 3458 98 3606 101
rect 3706 98 3798 101
rect 3810 98 3902 101
rect 4162 98 4358 101
rect 942 92 945 98
rect 530 88 550 91
rect 842 88 854 91
rect 858 88 942 91
rect 1026 88 1174 91
rect 1282 88 1342 91
rect 1362 88 1366 91
rect 1674 88 1790 91
rect 1882 88 2086 91
rect 2090 88 2121 91
rect 2194 88 2606 91
rect 2626 88 2670 91
rect 3070 91 3073 98
rect 2706 88 3073 91
rect 3346 88 3350 91
rect 3354 88 3534 91
rect 3570 88 3574 91
rect 3586 88 3590 91
rect 3610 88 3710 91
rect 3730 88 3966 91
rect 4202 88 4206 91
rect 354 78 358 81
rect 482 78 638 81
rect 922 78 998 81
rect 1002 78 1030 81
rect 1042 78 1118 81
rect 1230 81 1233 88
rect 1398 82 1401 88
rect 1230 78 1246 81
rect 1518 81 1521 88
rect 2118 82 2121 88
rect 2382 82 2385 88
rect 3078 82 3081 88
rect 1514 78 1521 81
rect 2050 78 2062 81
rect 2130 78 2150 81
rect 2154 78 2198 81
rect 2202 78 2302 81
rect 2402 78 2486 81
rect 2594 78 2606 81
rect 2634 78 2662 81
rect 2666 78 2670 81
rect 2682 78 2782 81
rect 2978 78 3006 81
rect 3214 81 3217 88
rect 4142 82 4145 88
rect 4150 82 4153 88
rect 3098 78 3217 81
rect 3226 78 3254 81
rect 3450 78 3638 81
rect 3650 78 3806 81
rect 3826 78 3902 81
rect 3962 78 4038 81
rect 4178 78 4246 81
rect 4250 78 4382 81
rect -26 71 -22 72
rect 30 71 33 78
rect -26 68 33 71
rect 158 72 161 78
rect 254 72 257 78
rect 1326 72 1329 78
rect 1502 72 1505 78
rect 346 68 374 71
rect 542 68 550 71
rect 634 68 806 71
rect 874 68 910 71
rect 978 68 1022 71
rect 1034 68 1086 71
rect 1106 68 1110 71
rect 1178 68 1302 71
rect 1378 68 1382 71
rect 1718 71 1721 78
rect 1718 68 1734 71
rect 1994 68 2014 71
rect 2170 68 2230 71
rect 2234 68 2238 71
rect 2258 68 2318 71
rect 2618 68 2694 71
rect 2698 68 2710 71
rect 2886 71 2889 78
rect 2758 68 2889 71
rect 2970 68 2974 71
rect 2994 68 3158 71
rect 3162 68 3198 71
rect 3218 68 3238 71
rect 3554 68 3614 71
rect 3682 68 3686 71
rect 3722 68 3726 71
rect 3882 68 4070 71
rect 4106 68 4166 71
rect 4186 68 4278 71
rect 4322 68 4326 71
rect 542 62 545 68
rect 2054 62 2057 68
rect 2758 62 2761 68
rect 374 58 382 61
rect 386 58 438 61
rect 586 58 678 61
rect 810 58 870 61
rect 874 58 934 61
rect 938 58 1014 61
rect 1018 58 1038 61
rect 1146 58 1270 61
rect 1314 58 1446 61
rect 1570 58 1662 61
rect 1778 58 1782 61
rect 1786 58 1830 61
rect 1898 58 1998 61
rect 2226 58 2278 61
rect 2282 58 2310 61
rect 2314 58 2342 61
rect 2346 58 2366 61
rect 2658 58 2678 61
rect 2786 58 2814 61
rect 2946 58 3038 61
rect 3170 58 3174 61
rect 3186 58 3238 61
rect 3338 58 3966 61
rect 3970 58 3998 61
rect 4122 58 4134 61
rect 4138 58 4206 61
rect 4314 58 4334 61
rect -26 51 -22 52
rect -26 48 6 51
rect 862 48 878 51
rect 1026 48 1030 51
rect 1066 48 1142 51
rect 1234 48 1598 51
rect 2010 48 2014 51
rect 2626 48 2638 51
rect 2662 48 2670 51
rect 2674 48 2742 51
rect 3274 48 3374 51
rect 3606 48 3614 51
rect 3618 48 3638 51
rect 3670 48 3694 51
rect 4162 48 4174 51
rect 862 42 865 48
rect 3670 42 3673 48
rect 1130 38 2022 41
rect 2026 38 2038 41
rect 2162 38 3190 41
rect 3194 38 3654 41
rect 4170 38 4174 41
rect 330 28 342 31
rect 1090 28 1326 31
rect 1346 28 2166 31
rect 2290 28 2294 31
rect 3234 28 3374 31
rect 1402 18 1414 21
rect 1434 18 2041 21
rect 2098 18 2310 21
rect 542 12 545 18
rect 558 12 561 18
rect 354 8 358 11
rect 434 8 446 11
rect 570 8 574 11
rect 634 8 638 11
rect 770 8 774 11
rect 1010 8 1014 11
rect 1194 8 1198 11
rect 1370 8 1374 11
rect 2038 11 2041 18
rect 2038 8 2134 11
rect 2154 8 2158 11
rect 2178 8 2398 11
rect 2506 8 2566 11
rect 2634 8 2638 11
rect 2746 8 2750 11
rect 4058 8 4070 11
rect 392 3 394 7
rect 398 3 401 7
rect 406 3 408 7
rect 1416 3 1418 7
rect 1422 3 1425 7
rect 1430 3 1432 7
rect 2440 3 2442 7
rect 2446 3 2449 7
rect 2454 3 2456 7
rect 3472 3 3474 7
rect 3478 3 3481 7
rect 3486 3 3488 7
<< m4contact >>
rect 898 3103 902 3107
rect 906 3103 909 3107
rect 909 3103 910 3107
rect 1930 3103 1934 3107
rect 1938 3103 1941 3107
rect 1941 3103 1942 3107
rect 2954 3103 2958 3107
rect 2962 3103 2965 3107
rect 2965 3103 2966 3107
rect 3978 3103 3982 3107
rect 3986 3103 3989 3107
rect 3989 3103 3990 3107
rect 1142 3098 1146 3102
rect 1174 3098 1178 3102
rect 1334 3098 1338 3102
rect 1702 3098 1706 3102
rect 1894 3098 1898 3102
rect 1910 3098 1914 3102
rect 2182 3098 2186 3102
rect 2502 3098 2506 3102
rect 2606 3098 2610 3102
rect 1470 3088 1474 3092
rect 2142 3088 2146 3092
rect 2406 3088 2410 3092
rect 4318 3088 4322 3092
rect 630 3078 634 3082
rect 4198 3078 4202 3082
rect 214 3068 218 3072
rect 550 3068 554 3072
rect 4166 3068 4170 3072
rect 4230 3068 4234 3072
rect 4246 3068 4250 3072
rect 4278 3068 4282 3072
rect 310 3058 314 3062
rect 710 3058 714 3062
rect 1598 3058 1602 3062
rect 1846 3058 1850 3062
rect 4158 3058 4162 3062
rect 3382 3048 3386 3052
rect 4030 3048 4034 3052
rect 4174 3048 4178 3052
rect 4262 3048 4266 3052
rect 4302 3048 4306 3052
rect 734 3038 738 3042
rect 3942 3038 3946 3042
rect 4182 3038 4186 3042
rect 1566 3028 1570 3032
rect 2278 3028 2282 3032
rect 4110 3028 4114 3032
rect 102 3018 106 3022
rect 1958 3018 1962 3022
rect 2470 3018 2474 3022
rect 3526 3018 3530 3022
rect 4262 3018 4266 3022
rect 4366 3018 4370 3022
rect 2926 3008 2930 3012
rect 394 3003 398 3007
rect 402 3003 405 3007
rect 405 3003 406 3007
rect 1418 3003 1422 3007
rect 1426 3003 1429 3007
rect 1429 3003 1430 3007
rect 2442 3003 2446 3007
rect 2450 3003 2453 3007
rect 2453 3003 2454 3007
rect 3474 3003 3478 3007
rect 3482 3003 3485 3007
rect 3485 3003 3486 3007
rect 2174 2998 2178 3002
rect 4142 2998 4146 3002
rect 4246 2998 4250 3002
rect 4302 2998 4306 3002
rect 3502 2988 3506 2992
rect 4094 2988 4098 2992
rect 2510 2978 2514 2982
rect 934 2968 938 2972
rect 1486 2968 1490 2972
rect 2046 2968 2050 2972
rect 2422 2968 2426 2972
rect 2806 2968 2810 2972
rect 4334 2968 4338 2972
rect 1462 2958 1466 2962
rect 2974 2958 2978 2962
rect 3742 2958 3746 2962
rect 3942 2958 3946 2962
rect 4134 2958 4138 2962
rect 4190 2958 4194 2962
rect 1670 2948 1674 2952
rect 2878 2948 2882 2952
rect 3070 2948 3074 2952
rect 3710 2948 3714 2952
rect 4150 2948 4154 2952
rect 4222 2948 4226 2952
rect 3342 2938 3346 2942
rect 702 2928 706 2932
rect 2166 2928 2170 2932
rect 2558 2928 2562 2932
rect 2758 2928 2762 2932
rect 2902 2928 2906 2932
rect 3390 2928 3394 2932
rect 3406 2928 3410 2932
rect 3694 2928 3698 2932
rect 3766 2928 3770 2932
rect 4214 2928 4218 2932
rect 4254 2928 4258 2932
rect 1246 2918 1250 2922
rect 1566 2918 1570 2922
rect 1878 2918 1882 2922
rect 2446 2918 2450 2922
rect 2750 2918 2754 2922
rect 3390 2918 3394 2922
rect 3726 2918 3730 2922
rect 1694 2908 1698 2912
rect 1830 2908 1834 2912
rect 2174 2908 2178 2912
rect 2318 2908 2322 2912
rect 2582 2908 2586 2912
rect 3542 2908 3546 2912
rect 3934 2908 3938 2912
rect 898 2903 902 2907
rect 906 2903 909 2907
rect 909 2903 910 2907
rect 1930 2903 1934 2907
rect 1938 2903 1941 2907
rect 1941 2903 1942 2907
rect 2954 2903 2958 2907
rect 2962 2903 2965 2907
rect 2965 2903 2966 2907
rect 3978 2903 3982 2907
rect 3986 2903 3989 2907
rect 3989 2903 3990 2907
rect 382 2898 386 2902
rect 2158 2898 2162 2902
rect 2414 2898 2418 2902
rect 2582 2898 2586 2902
rect 3598 2898 3602 2902
rect 934 2888 938 2892
rect 1478 2888 1482 2892
rect 2558 2888 2562 2892
rect 2886 2888 2890 2892
rect 3486 2888 3490 2892
rect 3582 2888 3586 2892
rect 3718 2888 3722 2892
rect 3550 2878 3554 2882
rect 3574 2878 3578 2882
rect 3638 2878 3642 2882
rect 3726 2878 3730 2882
rect 102 2868 106 2872
rect 878 2868 882 2872
rect 1198 2868 1202 2872
rect 1254 2868 1258 2872
rect 1750 2868 1754 2872
rect 3094 2868 3098 2872
rect 550 2858 554 2862
rect 1558 2858 1562 2862
rect 1886 2858 1890 2862
rect 2150 2858 2154 2862
rect 3350 2868 3354 2872
rect 3494 2868 3498 2872
rect 3918 2868 3922 2872
rect 4190 2868 4194 2872
rect 3526 2858 3530 2862
rect 3862 2858 3866 2862
rect 1022 2848 1026 2852
rect 1470 2848 1474 2852
rect 2462 2848 2466 2852
rect 2750 2848 2754 2852
rect 2758 2848 2762 2852
rect 4030 2848 4034 2852
rect 4270 2848 4274 2852
rect 534 2838 538 2842
rect 3254 2838 3258 2842
rect 3590 2838 3594 2842
rect 3942 2838 3946 2842
rect 2342 2828 2346 2832
rect 3550 2828 3554 2832
rect 3614 2828 3618 2832
rect 3638 2828 3642 2832
rect 726 2818 730 2822
rect 1270 2818 1274 2822
rect 1982 2818 1986 2822
rect 2670 2818 2674 2822
rect 3574 2818 3578 2822
rect 3654 2818 3658 2822
rect 3918 2818 3922 2822
rect 526 2808 530 2812
rect 1326 2808 1330 2812
rect 1438 2808 1442 2812
rect 1902 2808 1906 2812
rect 1998 2808 2002 2812
rect 3006 2808 3010 2812
rect 394 2803 398 2807
rect 402 2803 405 2807
rect 405 2803 406 2807
rect 1418 2803 1422 2807
rect 1426 2803 1429 2807
rect 1429 2803 1430 2807
rect 2442 2803 2446 2807
rect 2450 2803 2453 2807
rect 2453 2803 2454 2807
rect 3474 2803 3478 2807
rect 3482 2803 3485 2807
rect 3485 2803 3486 2807
rect 2062 2798 2066 2802
rect 4174 2798 4178 2802
rect 4358 2798 4362 2802
rect 30 2788 34 2792
rect 534 2788 538 2792
rect 1822 2788 1826 2792
rect 2246 2788 2250 2792
rect 2342 2788 2346 2792
rect 2910 2788 2914 2792
rect 3630 2788 3634 2792
rect 3798 2788 3802 2792
rect 4142 2788 4146 2792
rect 1918 2778 1922 2782
rect 3910 2778 3914 2782
rect 854 2768 858 2772
rect 1910 2768 1914 2772
rect 2094 2768 2098 2772
rect 2734 2768 2738 2772
rect 2806 2768 2810 2772
rect 3478 2768 3482 2772
rect 3790 2768 3794 2772
rect 4286 2768 4290 2772
rect 86 2758 90 2762
rect 214 2758 218 2762
rect 726 2758 730 2762
rect 1710 2758 1714 2762
rect 2462 2758 2466 2762
rect 4134 2758 4138 2762
rect 4238 2758 4242 2762
rect 4294 2758 4298 2762
rect 534 2748 538 2752
rect 758 2748 762 2752
rect 806 2748 810 2752
rect 886 2748 890 2752
rect 1014 2748 1018 2752
rect 2086 2748 2090 2752
rect 2110 2748 2114 2752
rect 2678 2748 2682 2752
rect 30 2738 34 2742
rect 2750 2748 2754 2752
rect 2822 2748 2826 2752
rect 3246 2748 3250 2752
rect 3542 2748 3546 2752
rect 3742 2748 3746 2752
rect 526 2738 530 2742
rect 574 2738 578 2742
rect 1166 2738 1170 2742
rect 1270 2738 1274 2742
rect 1622 2738 1626 2742
rect 1798 2738 1802 2742
rect 2054 2738 2058 2742
rect 2230 2738 2234 2742
rect 2566 2738 2570 2742
rect 2646 2738 2650 2742
rect 2742 2738 2746 2742
rect 2934 2738 2938 2742
rect 3094 2738 3098 2742
rect 3254 2738 3258 2742
rect 3502 2738 3506 2742
rect 3830 2738 3834 2742
rect 4062 2738 4066 2742
rect 4118 2738 4122 2742
rect 4246 2738 4250 2742
rect 4278 2738 4282 2742
rect 4334 2738 4338 2742
rect 422 2728 426 2732
rect 566 2728 570 2732
rect 1022 2728 1026 2732
rect 2150 2728 2154 2732
rect 2158 2728 2162 2732
rect 2318 2728 2322 2732
rect 2598 2728 2602 2732
rect 2942 2728 2946 2732
rect 2990 2728 2994 2732
rect 3198 2728 3202 2732
rect 3246 2728 3250 2732
rect 3422 2728 3426 2732
rect 3694 2728 3698 2732
rect 3726 2728 3730 2732
rect 3846 2728 3850 2732
rect 3958 2728 3962 2732
rect 4110 2728 4114 2732
rect 862 2718 866 2722
rect 1614 2718 1618 2722
rect 2918 2718 2922 2722
rect 3662 2718 3666 2722
rect 3702 2718 3706 2722
rect 3758 2718 3762 2722
rect 3966 2718 3970 2722
rect 4086 2718 4090 2722
rect 4094 2718 4098 2722
rect 4310 2718 4314 2722
rect 94 2708 98 2712
rect 1134 2708 1138 2712
rect 1254 2708 1258 2712
rect 1918 2708 1922 2712
rect 2398 2708 2402 2712
rect 2542 2708 2546 2712
rect 3998 2708 4002 2712
rect 4174 2708 4178 2712
rect 4206 2708 4210 2712
rect 4230 2708 4234 2712
rect 898 2703 902 2707
rect 906 2703 909 2707
rect 909 2703 910 2707
rect 1930 2703 1934 2707
rect 1938 2703 1941 2707
rect 1941 2703 1942 2707
rect 2954 2703 2958 2707
rect 2962 2703 2965 2707
rect 2965 2703 2966 2707
rect 3978 2703 3982 2707
rect 3986 2703 3989 2707
rect 3989 2703 3990 2707
rect 1046 2698 1050 2702
rect 1206 2698 1210 2702
rect 2630 2698 2634 2702
rect 2734 2698 2738 2702
rect 2998 2698 3002 2702
rect 3110 2698 3114 2702
rect 3998 2698 4002 2702
rect 4374 2698 4378 2702
rect 878 2688 882 2692
rect 886 2688 890 2692
rect 2222 2688 2226 2692
rect 2422 2688 2426 2692
rect 2590 2688 2594 2692
rect 4318 2688 4322 2692
rect 4382 2688 4386 2692
rect 4390 2688 4394 2692
rect 1398 2678 1402 2682
rect 1542 2678 1546 2682
rect 1766 2678 1770 2682
rect 2046 2678 2050 2682
rect 2054 2678 2058 2682
rect 2246 2678 2250 2682
rect 2654 2678 2658 2682
rect 3430 2678 3434 2682
rect 3614 2678 3618 2682
rect 3966 2678 3970 2682
rect 1238 2668 1242 2672
rect 1534 2668 1538 2672
rect 1662 2668 1666 2672
rect 1870 2668 1874 2672
rect 2414 2668 2418 2672
rect 2766 2668 2770 2672
rect 2942 2668 2946 2672
rect 3006 2668 3010 2672
rect 3062 2668 3066 2672
rect 4038 2668 4042 2672
rect 4206 2668 4210 2672
rect 534 2658 538 2662
rect 2230 2658 2234 2662
rect 2742 2658 2746 2662
rect 2750 2658 2754 2662
rect 2918 2658 2922 2662
rect 3158 2658 3162 2662
rect 3198 2658 3202 2662
rect 3742 2658 3746 2662
rect 518 2648 522 2652
rect 1182 2648 1186 2652
rect 1214 2648 1218 2652
rect 2350 2648 2354 2652
rect 2630 2648 2634 2652
rect 2790 2648 2794 2652
rect 3054 2648 3058 2652
rect 4102 2648 4106 2652
rect 4134 2648 4138 2652
rect 4150 2648 4154 2652
rect 4294 2648 4298 2652
rect 214 2638 218 2642
rect 574 2638 578 2642
rect 1302 2638 1306 2642
rect 2486 2638 2490 2642
rect 2742 2638 2746 2642
rect 2054 2628 2058 2632
rect 2254 2628 2258 2632
rect 2574 2628 2578 2632
rect 2814 2628 2818 2632
rect 3054 2628 3058 2632
rect 3126 2628 3130 2632
rect 3846 2628 3850 2632
rect 4190 2628 4194 2632
rect 1246 2618 1250 2622
rect 2182 2618 2186 2622
rect 2270 2618 2274 2622
rect 2750 2618 2754 2622
rect 2822 2618 2826 2622
rect 3774 2618 3778 2622
rect 3998 2618 4002 2622
rect 4086 2618 4090 2622
rect 1694 2608 1698 2612
rect 2406 2608 2410 2612
rect 2494 2608 2498 2612
rect 4022 2608 4026 2612
rect 4206 2608 4210 2612
rect 394 2603 398 2607
rect 402 2603 405 2607
rect 405 2603 406 2607
rect 1418 2603 1422 2607
rect 1426 2603 1429 2607
rect 1429 2603 1430 2607
rect 2442 2603 2446 2607
rect 2450 2603 2453 2607
rect 2453 2603 2454 2607
rect 3474 2603 3478 2607
rect 3482 2603 3485 2607
rect 3485 2603 3486 2607
rect 94 2598 98 2602
rect 606 2598 610 2602
rect 1190 2598 1194 2602
rect 2046 2598 2050 2602
rect 2238 2598 2242 2602
rect 2326 2598 2330 2602
rect 2974 2598 2978 2602
rect 3686 2598 3690 2602
rect 38 2588 42 2592
rect 1382 2588 1386 2592
rect 2070 2588 2074 2592
rect 2886 2588 2890 2592
rect 502 2578 506 2582
rect 590 2578 594 2582
rect 1542 2578 1546 2582
rect 2726 2578 2730 2582
rect 2822 2578 2826 2582
rect 3606 2578 3610 2582
rect 3854 2578 3858 2582
rect 4038 2578 4042 2582
rect 750 2568 754 2572
rect 1614 2568 1618 2572
rect 2214 2568 2218 2572
rect 2542 2568 2546 2572
rect 2630 2568 2634 2572
rect 4006 2568 4010 2572
rect 4134 2568 4138 2572
rect 110 2558 114 2562
rect 662 2558 666 2562
rect 1814 2558 1818 2562
rect 2014 2558 2018 2562
rect 2270 2558 2274 2562
rect 2502 2558 2506 2562
rect 2934 2558 2938 2562
rect 3254 2558 3258 2562
rect 3582 2558 3586 2562
rect 3718 2558 3722 2562
rect 3766 2558 3770 2562
rect 4310 2558 4314 2562
rect 4374 2558 4378 2562
rect 606 2548 610 2552
rect 758 2548 762 2552
rect 1750 2548 1754 2552
rect 1966 2548 1970 2552
rect 2646 2548 2650 2552
rect 2766 2548 2770 2552
rect 2806 2548 2810 2552
rect 3006 2548 3010 2552
rect 3230 2548 3234 2552
rect 3270 2548 3274 2552
rect 3598 2548 3602 2552
rect 4142 2548 4146 2552
rect 494 2538 498 2542
rect 510 2538 514 2542
rect 1134 2538 1138 2542
rect 1806 2538 1810 2542
rect 1918 2538 1922 2542
rect 1998 2538 2002 2542
rect 2062 2538 2066 2542
rect 2262 2538 2266 2542
rect 2326 2538 2330 2542
rect 2422 2538 2426 2542
rect 2542 2538 2546 2542
rect 2942 2538 2946 2542
rect 3718 2538 3722 2542
rect 3758 2538 3762 2542
rect 3838 2538 3842 2542
rect 4150 2538 4154 2542
rect 4310 2538 4314 2542
rect 486 2528 490 2532
rect 662 2528 666 2532
rect 1510 2528 1514 2532
rect 1630 2528 1634 2532
rect 1854 2528 1858 2532
rect 2094 2528 2098 2532
rect 2262 2528 2266 2532
rect 2294 2528 2298 2532
rect 2350 2528 2354 2532
rect 2422 2528 2426 2532
rect 2550 2528 2554 2532
rect 2598 2528 2602 2532
rect 2662 2528 2666 2532
rect 2974 2528 2978 2532
rect 3278 2528 3282 2532
rect 3390 2528 3394 2532
rect 3838 2528 3842 2532
rect 3894 2528 3898 2532
rect 4294 2528 4298 2532
rect 1550 2518 1554 2522
rect 2334 2518 2338 2522
rect 2598 2518 2602 2522
rect 2686 2518 2690 2522
rect 2694 2518 2698 2522
rect 3222 2518 3226 2522
rect 3502 2518 3506 2522
rect 3622 2518 3626 2522
rect 3854 2518 3858 2522
rect 574 2508 578 2512
rect 966 2508 970 2512
rect 2254 2508 2258 2512
rect 2478 2508 2482 2512
rect 2806 2508 2810 2512
rect 2942 2508 2946 2512
rect 3598 2508 3602 2512
rect 3790 2508 3794 2512
rect 3966 2508 3970 2512
rect 898 2503 902 2507
rect 906 2503 909 2507
rect 909 2503 910 2507
rect 1930 2503 1934 2507
rect 1938 2503 1941 2507
rect 1941 2503 1942 2507
rect 334 2498 338 2502
rect 1438 2498 1442 2502
rect 1446 2498 1450 2502
rect 2006 2498 2010 2502
rect 2954 2503 2958 2507
rect 2962 2503 2965 2507
rect 2965 2503 2966 2507
rect 3978 2503 3982 2507
rect 3986 2503 3989 2507
rect 3989 2503 3990 2507
rect 3846 2498 3850 2502
rect 582 2488 586 2492
rect 1230 2488 1234 2492
rect 1238 2488 1242 2492
rect 1622 2488 1626 2492
rect 1694 2488 1698 2492
rect 1734 2488 1738 2492
rect 1950 2488 1954 2492
rect 4190 2488 4194 2492
rect 86 2478 90 2482
rect 758 2478 762 2482
rect 1390 2478 1394 2482
rect 1686 2478 1690 2482
rect 2086 2478 2090 2482
rect 2638 2478 2642 2482
rect 3278 2478 3282 2482
rect 3534 2478 3538 2482
rect 3542 2478 3546 2482
rect 3910 2478 3914 2482
rect 4134 2478 4138 2482
rect 4238 2478 4242 2482
rect 1670 2468 1674 2472
rect 1854 2468 1858 2472
rect 1870 2468 1874 2472
rect 2518 2468 2522 2472
rect 2558 2468 2562 2472
rect 2702 2468 2706 2472
rect 2750 2468 2754 2472
rect 2998 2468 3002 2472
rect 3190 2468 3194 2472
rect 3198 2468 3202 2472
rect 3238 2468 3242 2472
rect 3326 2468 3330 2472
rect 3358 2468 3362 2472
rect 3694 2468 3698 2472
rect 4174 2468 4178 2472
rect 750 2458 754 2462
rect 1366 2458 1370 2462
rect 1662 2458 1666 2462
rect 1686 2458 1690 2462
rect 1838 2458 1842 2462
rect 2054 2458 2058 2462
rect 2118 2458 2122 2462
rect 2358 2458 2362 2462
rect 2366 2458 2370 2462
rect 2486 2458 2490 2462
rect 2782 2458 2786 2462
rect 2814 2458 2818 2462
rect 3246 2458 3250 2462
rect 3310 2458 3314 2462
rect 3318 2458 3322 2462
rect 3518 2458 3522 2462
rect 3534 2458 3538 2462
rect 3670 2458 3674 2462
rect 4174 2458 4178 2462
rect 38 2448 42 2452
rect 502 2448 506 2452
rect 622 2448 626 2452
rect 1070 2448 1074 2452
rect 1094 2448 1098 2452
rect 1350 2448 1354 2452
rect 1750 2448 1754 2452
rect 2078 2448 2082 2452
rect 2262 2448 2266 2452
rect 2334 2448 2338 2452
rect 2750 2448 2754 2452
rect 3062 2448 3066 2452
rect 3134 2448 3138 2452
rect 3190 2448 3194 2452
rect 4214 2448 4218 2452
rect 1654 2438 1658 2442
rect 1798 2438 1802 2442
rect 1902 2438 1906 2442
rect 2350 2438 2354 2442
rect 2798 2438 2802 2442
rect 2822 2438 2826 2442
rect 3270 2438 3274 2442
rect 590 2428 594 2432
rect 2110 2428 2114 2432
rect 2494 2428 2498 2432
rect 2758 2428 2762 2432
rect 3494 2428 3498 2432
rect 3662 2428 3666 2432
rect 3726 2428 3730 2432
rect 1830 2418 1834 2422
rect 2230 2418 2234 2422
rect 2310 2418 2314 2422
rect 3174 2418 3178 2422
rect 3406 2418 3410 2422
rect 3606 2418 3610 2422
rect 1510 2408 1514 2412
rect 1638 2408 1642 2412
rect 1998 2408 2002 2412
rect 2430 2408 2434 2412
rect 2646 2408 2650 2412
rect 2878 2408 2882 2412
rect 3310 2408 3314 2412
rect 3790 2408 3794 2412
rect 4262 2408 4266 2412
rect 394 2403 398 2407
rect 402 2403 405 2407
rect 405 2403 406 2407
rect 1418 2403 1422 2407
rect 1426 2403 1429 2407
rect 1429 2403 1430 2407
rect 1214 2398 1218 2402
rect 1398 2398 1402 2402
rect 2442 2403 2446 2407
rect 2450 2403 2453 2407
rect 2453 2403 2454 2407
rect 3474 2403 3478 2407
rect 3482 2403 3485 2407
rect 3485 2403 3486 2407
rect 1846 2398 1850 2402
rect 2422 2398 2426 2402
rect 2750 2398 2754 2402
rect 1406 2388 1410 2392
rect 1702 2388 1706 2392
rect 1950 2388 1954 2392
rect 2838 2388 2842 2392
rect 3734 2388 3738 2392
rect 4214 2388 4218 2392
rect 1134 2378 1138 2382
rect 1814 2378 1818 2382
rect 2062 2378 2066 2382
rect 2406 2378 2410 2382
rect 3014 2378 3018 2382
rect 3038 2378 3042 2382
rect 3614 2378 3618 2382
rect 4062 2378 4066 2382
rect 1142 2368 1146 2372
rect 1958 2368 1962 2372
rect 1974 2368 1978 2372
rect 2574 2368 2578 2372
rect 2646 2368 2650 2372
rect 2662 2368 2666 2372
rect 3254 2368 3258 2372
rect 3966 2368 3970 2372
rect 4358 2368 4362 2372
rect 1342 2358 1346 2362
rect 2486 2358 2490 2362
rect 2790 2358 2794 2362
rect 2974 2358 2978 2362
rect 3134 2358 3138 2362
rect 3166 2358 3170 2362
rect 4022 2358 4026 2362
rect 4374 2358 4378 2362
rect 1382 2348 1386 2352
rect 1686 2348 1690 2352
rect 1790 2348 1794 2352
rect 2078 2348 2082 2352
rect 2190 2348 2194 2352
rect 2326 2348 2330 2352
rect 2774 2348 2778 2352
rect 3086 2348 3090 2352
rect 3110 2348 3114 2352
rect 3902 2348 3906 2352
rect 4270 2348 4274 2352
rect 4382 2348 4386 2352
rect 174 2338 178 2342
rect 1062 2338 1066 2342
rect 1390 2338 1394 2342
rect 1398 2338 1402 2342
rect 1518 2338 1522 2342
rect 1630 2338 1634 2342
rect 1830 2338 1834 2342
rect 1862 2338 1866 2342
rect 1894 2338 1898 2342
rect 1990 2338 1994 2342
rect 2038 2338 2042 2342
rect 2094 2338 2098 2342
rect 2278 2338 2282 2342
rect 2462 2338 2466 2342
rect 2494 2338 2498 2342
rect 2630 2338 2634 2342
rect 2670 2338 2674 2342
rect 3078 2338 3082 2342
rect 3230 2338 3234 2342
rect 3358 2338 3362 2342
rect 3550 2338 3554 2342
rect 3566 2338 3570 2342
rect 3822 2338 3826 2342
rect 3870 2338 3874 2342
rect 4206 2338 4210 2342
rect 4318 2338 4322 2342
rect 86 2328 90 2332
rect 382 2328 386 2332
rect 574 2328 578 2332
rect 958 2328 962 2332
rect 1014 2328 1018 2332
rect 1142 2328 1146 2332
rect 1614 2328 1618 2332
rect 1622 2328 1626 2332
rect 1822 2328 1826 2332
rect 2086 2328 2090 2332
rect 2134 2328 2138 2332
rect 2230 2328 2234 2332
rect 2254 2328 2258 2332
rect 2342 2328 2346 2332
rect 2398 2328 2402 2332
rect 2678 2328 2682 2332
rect 2686 2328 2690 2332
rect 2822 2328 2826 2332
rect 3030 2328 3034 2332
rect 3182 2328 3186 2332
rect 3198 2328 3202 2332
rect 3686 2328 3690 2332
rect 3862 2328 3866 2332
rect 3894 2328 3898 2332
rect 4030 2328 4034 2332
rect 366 2318 370 2322
rect 726 2318 730 2322
rect 1158 2318 1162 2322
rect 1254 2318 1258 2322
rect 1662 2318 1666 2322
rect 2814 2318 2818 2322
rect 4038 2318 4042 2322
rect 4350 2318 4354 2322
rect 742 2308 746 2312
rect 1078 2308 1082 2312
rect 1670 2308 1674 2312
rect 1758 2308 1762 2312
rect 1846 2308 1850 2312
rect 1862 2308 1866 2312
rect 2134 2308 2138 2312
rect 2558 2308 2562 2312
rect 4254 2308 4258 2312
rect 4350 2308 4354 2312
rect 898 2303 902 2307
rect 906 2303 909 2307
rect 909 2303 910 2307
rect 1930 2303 1934 2307
rect 1938 2303 1941 2307
rect 1941 2303 1942 2307
rect 2954 2303 2958 2307
rect 2962 2303 2965 2307
rect 2965 2303 2966 2307
rect 3978 2303 3982 2307
rect 3986 2303 3989 2307
rect 3989 2303 3990 2307
rect 790 2298 794 2302
rect 1094 2298 1098 2302
rect 1438 2298 1442 2302
rect 1862 2298 1866 2302
rect 1982 2298 1986 2302
rect 2182 2298 2186 2302
rect 3702 2298 3706 2302
rect 3886 2298 3890 2302
rect 4062 2298 4066 2302
rect 1662 2288 1666 2292
rect 1678 2288 1682 2292
rect 3422 2288 3426 2292
rect 3430 2288 3434 2292
rect 4094 2288 4098 2292
rect 4166 2288 4170 2292
rect 166 2278 170 2282
rect 886 2278 890 2282
rect 950 2278 954 2282
rect 1022 2278 1026 2282
rect 1334 2278 1338 2282
rect 1646 2278 1650 2282
rect 1670 2278 1674 2282
rect 1694 2278 1698 2282
rect 1718 2278 1722 2282
rect 1774 2278 1778 2282
rect 2270 2278 2274 2282
rect 2502 2278 2506 2282
rect 2766 2278 2770 2282
rect 3854 2278 3858 2282
rect 3918 2278 3922 2282
rect 3990 2278 3994 2282
rect 4006 2278 4010 2282
rect 4206 2278 4210 2282
rect 4262 2278 4266 2282
rect 1198 2268 1202 2272
rect 1206 2268 1210 2272
rect 1302 2268 1306 2272
rect 1398 2268 1402 2272
rect 2222 2268 2226 2272
rect 2342 2268 2346 2272
rect 2398 2268 2402 2272
rect 3142 2268 3146 2272
rect 3550 2268 3554 2272
rect 3686 2268 3690 2272
rect 3742 2268 3746 2272
rect 4150 2268 4154 2272
rect 654 2258 658 2262
rect 798 2258 802 2262
rect 806 2258 810 2262
rect 830 2258 834 2262
rect 846 2258 850 2262
rect 1030 2258 1034 2262
rect 1126 2258 1130 2262
rect 1734 2258 1738 2262
rect 1870 2258 1874 2262
rect 2006 2258 2010 2262
rect 2014 2258 2018 2262
rect 2134 2258 2138 2262
rect 2374 2258 2378 2262
rect 2758 2258 2762 2262
rect 3006 2258 3010 2262
rect 3334 2258 3338 2262
rect 3350 2258 3354 2262
rect 3366 2258 3370 2262
rect 3398 2258 3402 2262
rect 4294 2258 4298 2262
rect 1310 2248 1314 2252
rect 1638 2248 1642 2252
rect 1686 2248 1690 2252
rect 1806 2248 1810 2252
rect 1982 2248 1986 2252
rect 2030 2248 2034 2252
rect 2198 2248 2202 2252
rect 3126 2248 3130 2252
rect 3302 2248 3306 2252
rect 854 2238 858 2242
rect 4062 2248 4066 2252
rect 1782 2238 1786 2242
rect 1902 2238 1906 2242
rect 2006 2238 2010 2242
rect 2014 2238 2018 2242
rect 2542 2238 2546 2242
rect 3606 2238 3610 2242
rect 590 2228 594 2232
rect 1310 2228 1314 2232
rect 1574 2228 1578 2232
rect 1774 2228 1778 2232
rect 1790 2228 1794 2232
rect 1990 2228 1994 2232
rect 2510 2228 2514 2232
rect 2750 2228 2754 2232
rect 2766 2228 2770 2232
rect 3198 2228 3202 2232
rect 3934 2228 3938 2232
rect 518 2218 522 2222
rect 974 2218 978 2222
rect 1014 2218 1018 2222
rect 1286 2218 1290 2222
rect 2406 2218 2410 2222
rect 2542 2218 2546 2222
rect 2846 2218 2850 2222
rect 4014 2218 4018 2222
rect 942 2208 946 2212
rect 1182 2208 1186 2212
rect 1358 2208 1362 2212
rect 1678 2208 1682 2212
rect 2286 2208 2290 2212
rect 3230 2208 3234 2212
rect 3238 2208 3242 2212
rect 3558 2208 3562 2212
rect 3846 2208 3850 2212
rect 394 2203 398 2207
rect 402 2203 405 2207
rect 405 2203 406 2207
rect 1418 2203 1422 2207
rect 1426 2203 1429 2207
rect 1429 2203 1430 2207
rect 2442 2203 2446 2207
rect 2450 2203 2453 2207
rect 2453 2203 2454 2207
rect 3474 2203 3478 2207
rect 3482 2203 3485 2207
rect 3485 2203 3486 2207
rect 422 2198 426 2202
rect 2006 2198 2010 2202
rect 2022 2198 2026 2202
rect 3430 2198 3434 2202
rect 3494 2198 3498 2202
rect 2318 2188 2322 2192
rect 2358 2188 2362 2192
rect 2878 2188 2882 2192
rect 3174 2188 3178 2192
rect 4022 2188 4026 2192
rect 702 2178 706 2182
rect 966 2178 970 2182
rect 1182 2178 1186 2182
rect 1622 2178 1626 2182
rect 2318 2178 2322 2182
rect 2366 2178 2370 2182
rect 3286 2178 3290 2182
rect 3774 2178 3778 2182
rect 846 2168 850 2172
rect 870 2168 874 2172
rect 1006 2168 1010 2172
rect 1054 2168 1058 2172
rect 2062 2168 2066 2172
rect 2118 2168 2122 2172
rect 2558 2168 2562 2172
rect 2998 2168 3002 2172
rect 4062 2168 4066 2172
rect 638 2158 642 2162
rect 1150 2158 1154 2162
rect 1438 2158 1442 2162
rect 1734 2158 1738 2162
rect 1766 2158 1770 2162
rect 2030 2158 2034 2162
rect 2150 2158 2154 2162
rect 2198 2158 2202 2162
rect 2406 2158 2410 2162
rect 2574 2158 2578 2162
rect 3158 2158 3162 2162
rect 3798 2158 3802 2162
rect 4070 2158 4074 2162
rect 22 2148 26 2152
rect 198 2148 202 2152
rect 814 2148 818 2152
rect 838 2148 842 2152
rect 862 2148 866 2152
rect 1382 2148 1386 2152
rect 182 2138 186 2142
rect 806 2138 810 2142
rect 878 2138 882 2142
rect 910 2138 914 2142
rect 918 2138 922 2142
rect 942 2138 946 2142
rect 1302 2138 1306 2142
rect 1902 2148 1906 2152
rect 2302 2148 2306 2152
rect 2670 2148 2674 2152
rect 2838 2148 2842 2152
rect 3206 2148 3210 2152
rect 3214 2148 3218 2152
rect 3294 2148 3298 2152
rect 3358 2148 3362 2152
rect 3542 2148 3546 2152
rect 3718 2148 3722 2152
rect 3774 2148 3778 2152
rect 3998 2148 4002 2152
rect 4054 2148 4058 2152
rect 4102 2148 4106 2152
rect 4366 2148 4370 2152
rect 2006 2138 2010 2142
rect 2254 2138 2258 2142
rect 2326 2138 2330 2142
rect 2582 2138 2586 2142
rect 2822 2138 2826 2142
rect 3710 2138 3714 2142
rect 3734 2138 3738 2142
rect 3966 2138 3970 2142
rect 174 2128 178 2132
rect 1166 2128 1170 2132
rect 1230 2128 1234 2132
rect 1526 2128 1530 2132
rect 1598 2128 1602 2132
rect 1998 2128 2002 2132
rect 2014 2128 2018 2132
rect 2062 2128 2066 2132
rect 2414 2128 2418 2132
rect 2558 2128 2562 2132
rect 2590 2128 2594 2132
rect 2790 2128 2794 2132
rect 2806 2128 2810 2132
rect 4078 2128 4082 2132
rect 4086 2128 4090 2132
rect 4222 2128 4226 2132
rect 4326 2128 4330 2132
rect 206 2118 210 2122
rect 494 2118 498 2122
rect 646 2118 650 2122
rect 654 2118 658 2122
rect 1174 2118 1178 2122
rect 1606 2118 1610 2122
rect 1702 2118 1706 2122
rect 2542 2118 2546 2122
rect 2654 2118 2658 2122
rect 582 2108 586 2112
rect 1062 2108 1066 2112
rect 1294 2108 1298 2112
rect 1534 2108 1538 2112
rect 1542 2108 1546 2112
rect 1910 2108 1914 2112
rect 2262 2108 2266 2112
rect 2326 2108 2330 2112
rect 2862 2108 2866 2112
rect 3310 2108 3314 2112
rect 3526 2108 3530 2112
rect 3958 2108 3962 2112
rect 898 2103 902 2107
rect 906 2103 909 2107
rect 909 2103 910 2107
rect 1930 2103 1934 2107
rect 1938 2103 1941 2107
rect 1941 2103 1942 2107
rect 2954 2103 2958 2107
rect 2962 2103 2965 2107
rect 2965 2103 2966 2107
rect 3978 2103 3982 2107
rect 3986 2103 3989 2107
rect 3989 2103 3990 2107
rect 1046 2098 1050 2102
rect 1518 2098 1522 2102
rect 1694 2098 1698 2102
rect 1886 2098 1890 2102
rect 1974 2098 1978 2102
rect 2214 2098 2218 2102
rect 2342 2098 2346 2102
rect 3134 2098 3138 2102
rect 4062 2098 4066 2102
rect 4166 2098 4170 2102
rect 4358 2098 4362 2102
rect 4374 2098 4378 2102
rect 1006 2088 1010 2092
rect 166 2078 170 2082
rect 646 2078 650 2082
rect 2110 2088 2114 2092
rect 2614 2088 2618 2092
rect 2710 2088 2714 2092
rect 2862 2088 2866 2092
rect 2886 2088 2890 2092
rect 3174 2088 3178 2092
rect 3190 2088 3194 2092
rect 3246 2088 3250 2092
rect 3254 2088 3258 2092
rect 3710 2088 3714 2092
rect 3822 2088 3826 2092
rect 4030 2088 4034 2092
rect 4062 2088 4066 2092
rect 934 2078 938 2082
rect 950 2078 954 2082
rect 1078 2078 1082 2082
rect 790 2068 794 2072
rect 798 2068 802 2072
rect 1710 2078 1714 2082
rect 1718 2078 1722 2082
rect 2302 2078 2306 2082
rect 2334 2078 2338 2082
rect 2374 2078 2378 2082
rect 2790 2078 2794 2082
rect 2822 2078 2826 2082
rect 3110 2078 3114 2082
rect 3238 2078 3242 2082
rect 3574 2078 3578 2082
rect 4110 2078 4114 2082
rect 4166 2078 4170 2082
rect 4222 2078 4226 2082
rect 4334 2078 4338 2082
rect 4366 2078 4370 2082
rect 1406 2068 1410 2072
rect 1470 2068 1474 2072
rect 1694 2068 1698 2072
rect 1726 2068 1730 2072
rect 2158 2068 2162 2072
rect 2446 2068 2450 2072
rect 2550 2068 2554 2072
rect 2686 2068 2690 2072
rect 2702 2068 2706 2072
rect 2758 2068 2762 2072
rect 3334 2068 3338 2072
rect 3510 2068 3514 2072
rect 3614 2068 3618 2072
rect 3646 2068 3650 2072
rect 3886 2068 3890 2072
rect 3950 2068 3954 2072
rect 3958 2068 3962 2072
rect 4006 2068 4010 2072
rect 4030 2068 4034 2072
rect 4046 2068 4050 2072
rect 4078 2068 4082 2072
rect 4326 2068 4330 2072
rect 534 2058 538 2062
rect 590 2058 594 2062
rect 750 2058 754 2062
rect 782 2058 786 2062
rect 1078 2058 1082 2062
rect 1286 2058 1290 2062
rect 1638 2058 1642 2062
rect 2086 2058 2090 2062
rect 2406 2058 2410 2062
rect 3814 2058 3818 2062
rect 3846 2058 3850 2062
rect 3886 2058 3890 2062
rect 4366 2058 4370 2062
rect 518 2048 522 2052
rect 678 2048 682 2052
rect 766 2048 770 2052
rect 878 2048 882 2052
rect 1166 2048 1170 2052
rect 1198 2048 1202 2052
rect 1822 2048 1826 2052
rect 1934 2048 1938 2052
rect 1966 2048 1970 2052
rect 2526 2048 2530 2052
rect 2766 2048 2770 2052
rect 2782 2048 2786 2052
rect 3238 2048 3242 2052
rect 3294 2048 3298 2052
rect 3350 2048 3354 2052
rect 3414 2048 3418 2052
rect 3462 2048 3466 2052
rect 3710 2048 3714 2052
rect 4062 2048 4066 2052
rect 982 2038 986 2042
rect 1174 2038 1178 2042
rect 1494 2038 1498 2042
rect 1518 2038 1522 2042
rect 1862 2038 1866 2042
rect 2662 2038 2666 2042
rect 2822 2038 2826 2042
rect 3798 2038 3802 2042
rect 4046 2038 4050 2042
rect 774 2028 778 2032
rect 934 2028 938 2032
rect 1014 2028 1018 2032
rect 1142 2028 1146 2032
rect 1902 2028 1906 2032
rect 2678 2028 2682 2032
rect 3126 2028 3130 2032
rect 3206 2028 3210 2032
rect 4014 2028 4018 2032
rect 4150 2028 4154 2032
rect 686 2018 690 2022
rect 814 2018 818 2022
rect 1118 2018 1122 2022
rect 2734 2018 2738 2022
rect 2750 2018 2754 2022
rect 2766 2018 2770 2022
rect 3094 2018 3098 2022
rect 638 2008 642 2012
rect 942 2008 946 2012
rect 1102 2008 1106 2012
rect 1838 2008 1842 2012
rect 1886 2008 1890 2012
rect 2030 2008 2034 2012
rect 2638 2008 2642 2012
rect 3462 2008 3466 2012
rect 3942 2008 3946 2012
rect 4238 2008 4242 2012
rect 394 2003 398 2007
rect 402 2003 405 2007
rect 405 2003 406 2007
rect 1418 2003 1422 2007
rect 1426 2003 1429 2007
rect 1429 2003 1430 2007
rect 2442 2003 2446 2007
rect 2450 2003 2453 2007
rect 2453 2003 2454 2007
rect 3474 2003 3478 2007
rect 3482 2003 3485 2007
rect 3485 2003 3486 2007
rect 6 1998 10 2002
rect 670 1998 674 2002
rect 702 1998 706 2002
rect 774 1998 778 2002
rect 1158 1998 1162 2002
rect 1558 1998 1562 2002
rect 1614 1998 1618 2002
rect 2174 1998 2178 2002
rect 2182 1998 2186 2002
rect 2630 1998 2634 2002
rect 3430 1998 3434 2002
rect 3590 1998 3594 2002
rect 774 1988 778 1992
rect 822 1988 826 1992
rect 1318 1988 1322 1992
rect 1750 1988 1754 1992
rect 1774 1988 1778 1992
rect 1854 1988 1858 1992
rect 1870 1988 1874 1992
rect 1942 1988 1946 1992
rect 990 1978 994 1982
rect 998 1978 1002 1982
rect 1454 1978 1458 1982
rect 1966 1978 1970 1982
rect 2158 1978 2162 1982
rect 2662 1978 2666 1982
rect 3646 1978 3650 1982
rect 670 1968 674 1972
rect 694 1968 698 1972
rect 718 1968 722 1972
rect 846 1968 850 1972
rect 1278 1968 1282 1972
rect 1310 1968 1314 1972
rect 1542 1968 1546 1972
rect 1606 1968 1610 1972
rect 2070 1968 2074 1972
rect 2574 1968 2578 1972
rect 2790 1968 2794 1972
rect 3094 1968 3098 1972
rect 3182 1968 3186 1972
rect 3342 1968 3346 1972
rect 3382 1968 3386 1972
rect 3766 1968 3770 1972
rect 4142 1968 4146 1972
rect 4166 1968 4170 1972
rect 4294 1968 4298 1972
rect 70 1958 74 1962
rect 726 1958 730 1962
rect 782 1958 786 1962
rect 1022 1958 1026 1962
rect 1142 1958 1146 1962
rect 1166 1958 1170 1962
rect 1574 1958 1578 1962
rect 2118 1958 2122 1962
rect 2638 1958 2642 1962
rect 2814 1958 2818 1962
rect 3086 1958 3090 1962
rect 3214 1958 3218 1962
rect 3606 1958 3610 1962
rect 3678 1958 3682 1962
rect 3950 1958 3954 1962
rect 4254 1958 4258 1962
rect 4310 1958 4314 1962
rect 6 1948 10 1952
rect 62 1948 66 1952
rect 174 1948 178 1952
rect 206 1948 210 1952
rect 718 1948 722 1952
rect 798 1948 802 1952
rect 806 1948 810 1952
rect 1366 1948 1370 1952
rect 1382 1948 1386 1952
rect 1750 1948 1754 1952
rect 1934 1948 1938 1952
rect 2038 1948 2042 1952
rect 2174 1948 2178 1952
rect 2590 1948 2594 1952
rect 2782 1948 2786 1952
rect 3150 1948 3154 1952
rect 3342 1948 3346 1952
rect 3718 1948 3722 1952
rect 4038 1948 4042 1952
rect 4094 1948 4098 1952
rect 4206 1948 4210 1952
rect 4342 1948 4346 1952
rect 166 1938 170 1942
rect 190 1938 194 1942
rect 926 1938 930 1942
rect 990 1938 994 1942
rect 1030 1938 1034 1942
rect 1134 1938 1138 1942
rect 1142 1938 1146 1942
rect 1158 1938 1162 1942
rect 1246 1938 1250 1942
rect 1270 1938 1274 1942
rect 1350 1938 1354 1942
rect 1366 1938 1370 1942
rect 1446 1938 1450 1942
rect 1734 1938 1738 1942
rect 1806 1938 1810 1942
rect 1910 1938 1914 1942
rect 1918 1938 1922 1942
rect 2014 1938 2018 1942
rect 2726 1938 2730 1942
rect 2902 1938 2906 1942
rect 2942 1938 2946 1942
rect 3182 1938 3186 1942
rect 3262 1938 3266 1942
rect 3318 1938 3322 1942
rect 3510 1938 3514 1942
rect 3614 1938 3618 1942
rect 3742 1938 3746 1942
rect 4078 1938 4082 1942
rect 4174 1938 4178 1942
rect 4254 1938 4258 1942
rect 334 1928 338 1932
rect 526 1928 530 1932
rect 710 1928 714 1932
rect 1302 1928 1306 1932
rect 1326 1928 1330 1932
rect 1438 1928 1442 1932
rect 1478 1928 1482 1932
rect 1582 1928 1586 1932
rect 1614 1928 1618 1932
rect 2166 1928 2170 1932
rect 2270 1928 2274 1932
rect 2278 1928 2282 1932
rect 2358 1928 2362 1932
rect 2430 1928 2434 1932
rect 2670 1928 2674 1932
rect 2806 1928 2810 1932
rect 3078 1928 3082 1932
rect 3150 1928 3154 1932
rect 3278 1928 3282 1932
rect 3542 1928 3546 1932
rect 3598 1928 3602 1932
rect 3798 1928 3802 1932
rect 3846 1928 3850 1932
rect 4262 1928 4266 1932
rect 822 1918 826 1922
rect 1758 1918 1762 1922
rect 2606 1918 2610 1922
rect 3750 1918 3754 1922
rect 4342 1918 4346 1922
rect 526 1908 530 1912
rect 598 1908 602 1912
rect 1110 1908 1114 1912
rect 1142 1908 1146 1912
rect 1382 1908 1386 1912
rect 1598 1908 1602 1912
rect 1654 1908 1658 1912
rect 1846 1908 1850 1912
rect 1918 1908 1922 1912
rect 2078 1908 2082 1912
rect 2382 1908 2386 1912
rect 2814 1908 2818 1912
rect 3166 1908 3170 1912
rect 3454 1908 3458 1912
rect 3878 1908 3882 1912
rect 3910 1908 3914 1912
rect 4062 1908 4066 1912
rect 898 1903 902 1907
rect 906 1903 909 1907
rect 909 1903 910 1907
rect 1930 1903 1934 1907
rect 1938 1903 1941 1907
rect 1941 1903 1942 1907
rect 2954 1903 2958 1907
rect 2962 1903 2965 1907
rect 2965 1903 2966 1907
rect 3978 1903 3982 1907
rect 3986 1903 3989 1907
rect 3989 1903 3990 1907
rect 534 1898 538 1902
rect 870 1898 874 1902
rect 1462 1898 1466 1902
rect 1614 1898 1618 1902
rect 1902 1898 1906 1902
rect 2430 1898 2434 1902
rect 2774 1898 2778 1902
rect 3222 1898 3226 1902
rect 3334 1898 3338 1902
rect 3494 1898 3498 1902
rect 4222 1898 4226 1902
rect 286 1888 290 1892
rect 1470 1888 1474 1892
rect 1566 1888 1570 1892
rect 3518 1888 3522 1892
rect 3526 1888 3530 1892
rect 3710 1888 3714 1892
rect 3734 1888 3738 1892
rect 3886 1888 3890 1892
rect 3910 1888 3914 1892
rect 4294 1888 4298 1892
rect 550 1878 554 1882
rect 1030 1878 1034 1882
rect 1126 1878 1130 1882
rect 1134 1878 1138 1882
rect 1318 1878 1322 1882
rect 1510 1878 1514 1882
rect 1526 1878 1530 1882
rect 1630 1878 1634 1882
rect 1766 1878 1770 1882
rect 1878 1878 1882 1882
rect 1918 1878 1922 1882
rect 2086 1878 2090 1882
rect 2126 1878 2130 1882
rect 2478 1878 2482 1882
rect 2518 1878 2522 1882
rect 2926 1878 2930 1882
rect 2974 1878 2978 1882
rect 190 1868 194 1872
rect 382 1868 386 1872
rect 534 1868 538 1872
rect 774 1868 778 1872
rect 838 1868 842 1872
rect 870 1868 874 1872
rect 1006 1868 1010 1872
rect 1726 1868 1730 1872
rect 726 1858 730 1862
rect 782 1858 786 1862
rect 1006 1858 1010 1862
rect 1070 1858 1074 1862
rect 1206 1858 1210 1862
rect 1286 1858 1290 1862
rect 1294 1858 1298 1862
rect 1462 1858 1466 1862
rect 2366 1868 2370 1872
rect 2790 1868 2794 1872
rect 3494 1878 3498 1882
rect 3798 1878 3802 1882
rect 3814 1878 3818 1882
rect 4142 1878 4146 1882
rect 4166 1878 4170 1882
rect 3526 1868 3530 1872
rect 3726 1868 3730 1872
rect 3798 1868 3802 1872
rect 4326 1868 4330 1872
rect 1694 1858 1698 1862
rect 1750 1858 1754 1862
rect 2006 1858 2010 1862
rect 2070 1858 2074 1862
rect 2470 1858 2474 1862
rect 3622 1858 3626 1862
rect 3734 1858 3738 1862
rect 3750 1858 3754 1862
rect 4102 1858 4106 1862
rect 550 1848 554 1852
rect 1470 1848 1474 1852
rect 1534 1848 1538 1852
rect 1662 1848 1666 1852
rect 2054 1848 2058 1852
rect 2094 1848 2098 1852
rect 2102 1848 2106 1852
rect 2246 1848 2250 1852
rect 2462 1848 2466 1852
rect 3654 1848 3658 1852
rect 3830 1848 3834 1852
rect 4238 1848 4242 1852
rect 790 1838 794 1842
rect 1374 1838 1378 1842
rect 1414 1838 1418 1842
rect 1454 1838 1458 1842
rect 1478 1838 1482 1842
rect 1638 1838 1642 1842
rect 2646 1838 2650 1842
rect 2654 1838 2658 1842
rect 3014 1838 3018 1842
rect 3918 1838 3922 1842
rect 918 1828 922 1832
rect 1342 1828 1346 1832
rect 3694 1828 3698 1832
rect 3702 1828 3706 1832
rect 798 1818 802 1822
rect 1318 1818 1322 1822
rect 1342 1818 1346 1822
rect 1854 1818 1858 1822
rect 2070 1818 2074 1822
rect 2510 1818 2514 1822
rect 3054 1818 3058 1822
rect 3406 1818 3410 1822
rect 3710 1818 3714 1822
rect 3750 1818 3754 1822
rect 686 1808 690 1812
rect 1230 1808 1234 1812
rect 1894 1808 1898 1812
rect 2102 1808 2106 1812
rect 2654 1808 2658 1812
rect 3526 1808 3530 1812
rect 394 1803 398 1807
rect 402 1803 405 1807
rect 405 1803 406 1807
rect 1418 1803 1422 1807
rect 1426 1803 1429 1807
rect 1429 1803 1430 1807
rect 2442 1803 2446 1807
rect 2450 1803 2453 1807
rect 2453 1803 2454 1807
rect 3474 1803 3478 1807
rect 3482 1803 3485 1807
rect 3485 1803 3486 1807
rect 1270 1798 1274 1802
rect 1350 1798 1354 1802
rect 1686 1798 1690 1802
rect 2166 1798 2170 1802
rect 2406 1798 2410 1802
rect 2462 1798 2466 1802
rect 3062 1798 3066 1802
rect 3190 1798 3194 1802
rect 3598 1798 3602 1802
rect 4038 1798 4042 1802
rect 4150 1798 4154 1802
rect 6 1788 10 1792
rect 702 1788 706 1792
rect 1206 1788 1210 1792
rect 2518 1788 2522 1792
rect 2646 1788 2650 1792
rect 3742 1788 3746 1792
rect 854 1778 858 1782
rect 1774 1778 1778 1782
rect 2054 1778 2058 1782
rect 2190 1778 2194 1782
rect 2318 1778 2322 1782
rect 3422 1778 3426 1782
rect 3734 1778 3738 1782
rect 4294 1778 4298 1782
rect 4358 1778 4362 1782
rect 734 1768 738 1772
rect 982 1768 986 1772
rect 1838 1768 1842 1772
rect 1854 1768 1858 1772
rect 2078 1768 2082 1772
rect 2150 1768 2154 1772
rect 2182 1768 2186 1772
rect 3750 1768 3754 1772
rect 3782 1768 3786 1772
rect 4046 1768 4050 1772
rect 4086 1768 4090 1772
rect 974 1758 978 1762
rect 1070 1758 1074 1762
rect 1126 1758 1130 1762
rect 1158 1758 1162 1762
rect 1486 1758 1490 1762
rect 1510 1758 1514 1762
rect 1662 1758 1666 1762
rect 1990 1758 1994 1762
rect 2046 1758 2050 1762
rect 2230 1758 2234 1762
rect 2246 1758 2250 1762
rect 2454 1758 2458 1762
rect 2590 1758 2594 1762
rect 2702 1758 2706 1762
rect 2766 1758 2770 1762
rect 3094 1758 3098 1762
rect 3294 1758 3298 1762
rect 3790 1758 3794 1762
rect 4110 1758 4114 1762
rect 4174 1758 4178 1762
rect 886 1748 890 1752
rect 1326 1748 1330 1752
rect 1374 1748 1378 1752
rect 1486 1748 1490 1752
rect 1662 1748 1666 1752
rect 2054 1748 2058 1752
rect 2150 1748 2154 1752
rect 2902 1748 2906 1752
rect 3118 1748 3122 1752
rect 3654 1748 3658 1752
rect 3670 1748 3674 1752
rect 3774 1748 3778 1752
rect 4246 1748 4250 1752
rect 4390 1748 4394 1752
rect 158 1738 162 1742
rect 750 1738 754 1742
rect 1046 1738 1050 1742
rect 1974 1738 1978 1742
rect 2102 1738 2106 1742
rect 2166 1738 2170 1742
rect 2190 1738 2194 1742
rect 2254 1738 2258 1742
rect 2350 1738 2354 1742
rect 2750 1738 2754 1742
rect 3182 1738 3186 1742
rect 3614 1738 3618 1742
rect 3726 1738 3730 1742
rect 3766 1738 3770 1742
rect 4102 1738 4106 1742
rect 574 1728 578 1732
rect 718 1728 722 1732
rect 806 1728 810 1732
rect 902 1728 906 1732
rect 966 1728 970 1732
rect 1014 1728 1018 1732
rect 1062 1728 1066 1732
rect 1070 1728 1074 1732
rect 1246 1728 1250 1732
rect 1366 1728 1370 1732
rect 1526 1728 1530 1732
rect 1582 1728 1586 1732
rect 1702 1728 1706 1732
rect 1846 1728 1850 1732
rect 1958 1728 1962 1732
rect 1982 1728 1986 1732
rect 2006 1728 2010 1732
rect 2686 1728 2690 1732
rect 3126 1728 3130 1732
rect 3278 1728 3282 1732
rect 3590 1728 3594 1732
rect 3702 1728 3706 1732
rect 4046 1728 4050 1732
rect 4198 1728 4202 1732
rect 526 1718 530 1722
rect 926 1718 930 1722
rect 950 1718 954 1722
rect 966 1718 970 1722
rect 1022 1718 1026 1722
rect 1166 1718 1170 1722
rect 1390 1718 1394 1722
rect 1534 1718 1538 1722
rect 1678 1718 1682 1722
rect 1790 1718 1794 1722
rect 1806 1718 1810 1722
rect 2366 1718 2370 1722
rect 3102 1718 3106 1722
rect 3430 1718 3434 1722
rect 3446 1718 3450 1722
rect 4302 1718 4306 1722
rect 1574 1708 1578 1712
rect 2990 1708 2994 1712
rect 3414 1708 3418 1712
rect 3678 1708 3682 1712
rect 3902 1708 3906 1712
rect 898 1703 902 1707
rect 906 1703 909 1707
rect 909 1703 910 1707
rect 1930 1703 1934 1707
rect 1938 1703 1941 1707
rect 1941 1703 1942 1707
rect 790 1688 794 1692
rect 1334 1698 1338 1702
rect 1654 1698 1658 1702
rect 1886 1698 1890 1702
rect 2006 1698 2010 1702
rect 2046 1698 2050 1702
rect 2174 1698 2178 1702
rect 2238 1698 2242 1702
rect 2954 1703 2958 1707
rect 2962 1703 2965 1707
rect 2965 1703 2966 1707
rect 2710 1698 2714 1702
rect 3302 1698 3306 1702
rect 3510 1698 3514 1702
rect 3978 1703 3982 1707
rect 3986 1703 3989 1707
rect 3989 1703 3990 1707
rect 4358 1698 4362 1702
rect 982 1688 986 1692
rect 1134 1688 1138 1692
rect 1790 1688 1794 1692
rect 1806 1688 1810 1692
rect 1926 1688 1930 1692
rect 2254 1688 2258 1692
rect 2278 1688 2282 1692
rect 2742 1688 2746 1692
rect 2774 1688 2778 1692
rect 3454 1688 3458 1692
rect 3502 1688 3506 1692
rect 3822 1688 3826 1692
rect 166 1678 170 1682
rect 718 1678 722 1682
rect 766 1678 770 1682
rect 1102 1678 1106 1682
rect 1206 1678 1210 1682
rect 1286 1678 1290 1682
rect 1302 1678 1306 1682
rect 1318 1678 1322 1682
rect 1446 1678 1450 1682
rect 1654 1678 1658 1682
rect 2014 1678 2018 1682
rect 2646 1678 2650 1682
rect 2926 1678 2930 1682
rect 3166 1678 3170 1682
rect 3478 1678 3482 1682
rect 3622 1678 3626 1682
rect 3750 1678 3754 1682
rect 3926 1678 3930 1682
rect 4246 1678 4250 1682
rect 158 1668 162 1672
rect 582 1668 586 1672
rect 606 1668 610 1672
rect 734 1668 738 1672
rect 1014 1668 1018 1672
rect 1142 1668 1146 1672
rect 1366 1668 1370 1672
rect 1438 1668 1442 1672
rect 1526 1668 1530 1672
rect 1686 1668 1690 1672
rect 1702 1668 1706 1672
rect 2262 1668 2266 1672
rect 2582 1668 2586 1672
rect 4110 1668 4114 1672
rect 4262 1668 4266 1672
rect 166 1658 170 1662
rect 630 1658 634 1662
rect 814 1658 818 1662
rect 910 1658 914 1662
rect 934 1658 938 1662
rect 958 1658 962 1662
rect 1374 1658 1378 1662
rect 1382 1658 1386 1662
rect 1454 1658 1458 1662
rect 1510 1658 1514 1662
rect 1606 1658 1610 1662
rect 1694 1658 1698 1662
rect 2038 1658 2042 1662
rect 2102 1658 2106 1662
rect 2654 1658 2658 1662
rect 3150 1658 3154 1662
rect 3214 1658 3218 1662
rect 3270 1658 3274 1662
rect 3422 1658 3426 1662
rect 3638 1658 3642 1662
rect 6 1648 10 1652
rect 646 1648 650 1652
rect 878 1648 882 1652
rect 974 1648 978 1652
rect 1102 1648 1106 1652
rect 1126 1648 1130 1652
rect 1214 1648 1218 1652
rect 1366 1648 1370 1652
rect 1494 1648 1498 1652
rect 1774 1648 1778 1652
rect 1782 1648 1786 1652
rect 1910 1648 1914 1652
rect 2006 1648 2010 1652
rect 2374 1648 2378 1652
rect 2718 1648 2722 1652
rect 2830 1648 2834 1652
rect 2870 1648 2874 1652
rect 3182 1648 3186 1652
rect 3470 1648 3474 1652
rect 3598 1648 3602 1652
rect 3686 1648 3690 1652
rect 3950 1648 3954 1652
rect 4030 1648 4034 1652
rect 4046 1648 4050 1652
rect 4126 1648 4130 1652
rect 4142 1648 4146 1652
rect 4286 1648 4290 1652
rect 4366 1648 4370 1652
rect 710 1638 714 1642
rect 1190 1638 1194 1642
rect 1406 1638 1410 1642
rect 1462 1638 1466 1642
rect 1758 1638 1762 1642
rect 1862 1638 1866 1642
rect 2110 1638 2114 1642
rect 2134 1638 2138 1642
rect 2590 1638 2594 1642
rect 2790 1638 2794 1642
rect 3246 1638 3250 1642
rect 3502 1638 3506 1642
rect 4366 1638 4370 1642
rect 838 1628 842 1632
rect 870 1628 874 1632
rect 1262 1628 1266 1632
rect 1534 1628 1538 1632
rect 1582 1628 1586 1632
rect 1966 1628 1970 1632
rect 2198 1628 2202 1632
rect 2222 1628 2226 1632
rect 3086 1628 3090 1632
rect 4310 1628 4314 1632
rect 4358 1628 4362 1632
rect 6 1618 10 1622
rect 1814 1618 1818 1622
rect 1838 1618 1842 1622
rect 1918 1618 1922 1622
rect 1966 1618 1970 1622
rect 2070 1618 2074 1622
rect 2598 1618 2602 1622
rect 2910 1618 2914 1622
rect 2974 1618 2978 1622
rect 3126 1618 3130 1622
rect 4302 1618 4306 1622
rect 1406 1608 1410 1612
rect 2086 1608 2090 1612
rect 2118 1608 2122 1612
rect 2566 1608 2570 1612
rect 3134 1608 3138 1612
rect 4310 1608 4314 1612
rect 394 1603 398 1607
rect 402 1603 405 1607
rect 405 1603 406 1607
rect 1418 1603 1422 1607
rect 1426 1603 1429 1607
rect 1429 1603 1430 1607
rect 2442 1603 2446 1607
rect 2450 1603 2453 1607
rect 2453 1603 2454 1607
rect 3474 1603 3478 1607
rect 3482 1603 3485 1607
rect 3485 1603 3486 1607
rect 774 1598 778 1602
rect 1462 1598 1466 1602
rect 1542 1598 1546 1602
rect 1638 1598 1642 1602
rect 1654 1598 1658 1602
rect 1990 1598 1994 1602
rect 2182 1598 2186 1602
rect 2422 1598 2426 1602
rect 2878 1598 2882 1602
rect 2886 1598 2890 1602
rect 854 1588 858 1592
rect 1086 1588 1090 1592
rect 1118 1588 1122 1592
rect 1406 1588 1410 1592
rect 1646 1588 1650 1592
rect 1662 1588 1666 1592
rect 3126 1588 3130 1592
rect 3822 1588 3826 1592
rect 4286 1588 4290 1592
rect 4326 1588 4330 1592
rect 950 1578 954 1582
rect 1494 1578 1498 1582
rect 2878 1578 2882 1582
rect 3462 1578 3466 1582
rect 766 1568 770 1572
rect 798 1568 802 1572
rect 806 1568 810 1572
rect 838 1568 842 1572
rect 1630 1568 1634 1572
rect 1718 1568 1722 1572
rect 3166 1568 3170 1572
rect 3294 1568 3298 1572
rect 3702 1568 3706 1572
rect 3886 1568 3890 1572
rect 4326 1568 4330 1572
rect 430 1558 434 1562
rect 1358 1558 1362 1562
rect 1502 1558 1506 1562
rect 1734 1558 1738 1562
rect 1998 1558 2002 1562
rect 2150 1558 2154 1562
rect 2198 1558 2202 1562
rect 2302 1558 2306 1562
rect 2822 1558 2826 1562
rect 2838 1558 2842 1562
rect 3206 1558 3210 1562
rect 3310 1558 3314 1562
rect 3334 1558 3338 1562
rect 3838 1558 3842 1562
rect 3934 1558 3938 1562
rect 4046 1558 4050 1562
rect 4190 1558 4194 1562
rect 14 1548 18 1552
rect 174 1548 178 1552
rect 862 1548 866 1552
rect 902 1548 906 1552
rect 1462 1548 1466 1552
rect 1510 1548 1514 1552
rect 1550 1548 1554 1552
rect 1654 1548 1658 1552
rect 1662 1548 1666 1552
rect 1814 1548 1818 1552
rect 1894 1548 1898 1552
rect 2582 1548 2586 1552
rect 2622 1548 2626 1552
rect 2718 1548 2722 1552
rect 2894 1548 2898 1552
rect 3326 1548 3330 1552
rect 3398 1548 3402 1552
rect 3414 1548 3418 1552
rect 3550 1548 3554 1552
rect 3574 1548 3578 1552
rect 3638 1548 3642 1552
rect 3838 1548 3842 1552
rect 4246 1548 4250 1552
rect 102 1538 106 1542
rect 614 1538 618 1542
rect 686 1538 690 1542
rect 718 1538 722 1542
rect 838 1538 842 1542
rect 926 1538 930 1542
rect 1262 1538 1266 1542
rect 1438 1538 1442 1542
rect 1446 1538 1450 1542
rect 1478 1538 1482 1542
rect 1678 1538 1682 1542
rect 1798 1538 1802 1542
rect 1830 1538 1834 1542
rect 1838 1538 1842 1542
rect 1926 1538 1930 1542
rect 1958 1538 1962 1542
rect 2094 1538 2098 1542
rect 2366 1538 2370 1542
rect 2470 1538 2474 1542
rect 3070 1538 3074 1542
rect 3582 1538 3586 1542
rect 3622 1538 3626 1542
rect 3758 1538 3762 1542
rect 3926 1538 3930 1542
rect 4166 1538 4170 1542
rect 198 1528 202 1532
rect 574 1528 578 1532
rect 638 1528 642 1532
rect 1134 1528 1138 1532
rect 1582 1528 1586 1532
rect 1990 1528 1994 1532
rect 2206 1528 2210 1532
rect 2422 1528 2426 1532
rect 2598 1528 2602 1532
rect 2790 1528 2794 1532
rect 3054 1528 3058 1532
rect 3142 1528 3146 1532
rect 3166 1528 3170 1532
rect 3190 1528 3194 1532
rect 3198 1528 3202 1532
rect 3318 1528 3322 1532
rect 3342 1528 3346 1532
rect 3350 1528 3354 1532
rect 3358 1528 3362 1532
rect 3502 1528 3506 1532
rect 3510 1528 3514 1532
rect 3534 1528 3538 1532
rect 3590 1528 3594 1532
rect 3622 1528 3626 1532
rect 3686 1528 3690 1532
rect 422 1518 426 1522
rect 838 1518 842 1522
rect 1078 1518 1082 1522
rect 1238 1518 1242 1522
rect 1606 1518 1610 1522
rect 1974 1518 1978 1522
rect 2342 1518 2346 1522
rect 2558 1518 2562 1522
rect 2846 1518 2850 1522
rect 2942 1518 2946 1522
rect 3166 1518 3170 1522
rect 3374 1518 3378 1522
rect 3414 1518 3418 1522
rect 3502 1518 3506 1522
rect 3558 1518 3562 1522
rect 6 1508 10 1512
rect 1406 1508 1410 1512
rect 1622 1508 1626 1512
rect 1686 1508 1690 1512
rect 1726 1508 1730 1512
rect 1790 1508 1794 1512
rect 1910 1508 1914 1512
rect 1974 1508 1978 1512
rect 2302 1508 2306 1512
rect 3462 1508 3466 1512
rect 3478 1508 3482 1512
rect 3614 1508 3618 1512
rect 3742 1508 3746 1512
rect 898 1503 902 1507
rect 906 1503 909 1507
rect 909 1503 910 1507
rect 1930 1503 1934 1507
rect 1938 1503 1941 1507
rect 1941 1503 1942 1507
rect 2954 1503 2958 1507
rect 2962 1503 2965 1507
rect 2965 1503 2966 1507
rect 3978 1503 3982 1507
rect 3986 1503 3989 1507
rect 3989 1503 3990 1507
rect 614 1498 618 1502
rect 814 1498 818 1502
rect 838 1498 842 1502
rect 886 1498 890 1502
rect 982 1498 986 1502
rect 1462 1498 1466 1502
rect 1622 1498 1626 1502
rect 2246 1498 2250 1502
rect 2974 1498 2978 1502
rect 6 1488 10 1492
rect 14 1488 18 1492
rect 1190 1488 1194 1492
rect 1390 1488 1394 1492
rect 1678 1488 1682 1492
rect 1782 1488 1786 1492
rect 2382 1488 2386 1492
rect 2558 1488 2562 1492
rect 2606 1488 2610 1492
rect 2814 1488 2818 1492
rect 2982 1488 2986 1492
rect 3550 1488 3554 1492
rect 3710 1488 3714 1492
rect 3734 1488 3738 1492
rect 830 1478 834 1482
rect 1518 1478 1522 1482
rect 1534 1478 1538 1482
rect 1710 1478 1714 1482
rect 1758 1478 1762 1482
rect 1886 1478 1890 1482
rect 2190 1478 2194 1482
rect 54 1468 58 1472
rect 166 1468 170 1472
rect 2830 1478 2834 1482
rect 3278 1478 3282 1482
rect 3318 1478 3322 1482
rect 3358 1478 3362 1482
rect 3678 1478 3682 1482
rect 3830 1478 3834 1482
rect 3942 1478 3946 1482
rect 4134 1478 4138 1482
rect 4198 1478 4202 1482
rect 4214 1478 4218 1482
rect 414 1468 418 1472
rect 654 1468 658 1472
rect 750 1468 754 1472
rect 1366 1468 1370 1472
rect 1494 1468 1498 1472
rect 1774 1468 1778 1472
rect 1894 1468 1898 1472
rect 2406 1468 2410 1472
rect 2830 1468 2834 1472
rect 3030 1468 3034 1472
rect 3110 1468 3114 1472
rect 3222 1468 3226 1472
rect 3302 1468 3306 1472
rect 3334 1468 3338 1472
rect 3366 1468 3370 1472
rect 3406 1468 3410 1472
rect 3430 1468 3434 1472
rect 3806 1468 3810 1472
rect 4270 1468 4274 1472
rect 4302 1468 4306 1472
rect 510 1458 514 1462
rect 598 1458 602 1462
rect 622 1458 626 1462
rect 726 1458 730 1462
rect 774 1458 778 1462
rect 958 1458 962 1462
rect 1142 1458 1146 1462
rect 1254 1458 1258 1462
rect 1406 1458 1410 1462
rect 1566 1458 1570 1462
rect 1590 1458 1594 1462
rect 1686 1458 1690 1462
rect 1942 1458 1946 1462
rect 2390 1458 2394 1462
rect 2718 1458 2722 1462
rect 2726 1458 2730 1462
rect 2822 1458 2826 1462
rect 2870 1458 2874 1462
rect 2902 1458 2906 1462
rect 4086 1458 4090 1462
rect 4230 1458 4234 1462
rect 4238 1458 4242 1462
rect 4302 1458 4306 1462
rect 78 1448 82 1452
rect 606 1448 610 1452
rect 1454 1448 1458 1452
rect 1470 1448 1474 1452
rect 1646 1448 1650 1452
rect 1662 1448 1666 1452
rect 1782 1448 1786 1452
rect 1790 1448 1794 1452
rect 2006 1448 2010 1452
rect 2414 1448 2418 1452
rect 3318 1448 3322 1452
rect 3334 1448 3338 1452
rect 3358 1448 3362 1452
rect 3950 1448 3954 1452
rect 518 1438 522 1442
rect 550 1438 554 1442
rect 790 1438 794 1442
rect 1406 1438 1410 1442
rect 1502 1438 1506 1442
rect 1670 1438 1674 1442
rect 1870 1438 1874 1442
rect 1910 1438 1914 1442
rect 1990 1438 1994 1442
rect 2494 1438 2498 1442
rect 3414 1438 3418 1442
rect 3630 1438 3634 1442
rect 3646 1438 3650 1442
rect 3758 1438 3762 1442
rect 3910 1438 3914 1442
rect 710 1428 714 1432
rect 2886 1428 2890 1432
rect 3598 1428 3602 1432
rect 694 1418 698 1422
rect 886 1418 890 1422
rect 2526 1418 2530 1422
rect 2854 1418 2858 1422
rect 3374 1418 3378 1422
rect 3438 1418 3442 1422
rect 3622 1418 3626 1422
rect 4190 1418 4194 1422
rect 414 1408 418 1412
rect 1302 1408 1306 1412
rect 1438 1408 1442 1412
rect 2262 1408 2266 1412
rect 2590 1408 2594 1412
rect 2742 1408 2746 1412
rect 394 1403 398 1407
rect 402 1403 405 1407
rect 405 1403 406 1407
rect 1418 1403 1422 1407
rect 1426 1403 1429 1407
rect 1429 1403 1430 1407
rect 2442 1403 2446 1407
rect 2450 1403 2453 1407
rect 2453 1403 2454 1407
rect 870 1398 874 1402
rect 1470 1398 1474 1402
rect 3474 1403 3478 1407
rect 3482 1403 3485 1407
rect 3485 1403 3486 1407
rect 2934 1398 2938 1402
rect 2974 1398 2978 1402
rect 3094 1398 3098 1402
rect 3494 1398 3498 1402
rect 486 1388 490 1392
rect 1718 1388 1722 1392
rect 1750 1388 1754 1392
rect 1918 1388 1922 1392
rect 2006 1388 2010 1392
rect 2350 1388 2354 1392
rect 2382 1388 2386 1392
rect 2494 1388 2498 1392
rect 2838 1388 2842 1392
rect 2846 1388 2850 1392
rect 3390 1388 3394 1392
rect 1462 1378 1466 1382
rect 1494 1378 1498 1382
rect 1638 1378 1642 1382
rect 1646 1378 1650 1382
rect 1726 1378 1730 1382
rect 2102 1378 2106 1382
rect 2118 1378 2122 1382
rect 2486 1378 2490 1382
rect 4086 1378 4090 1382
rect 798 1368 802 1372
rect 1046 1368 1050 1372
rect 1222 1368 1226 1372
rect 2630 1368 2634 1372
rect 3030 1368 3034 1372
rect 3198 1368 3202 1372
rect 3526 1368 3530 1372
rect 4038 1368 4042 1372
rect 4054 1368 4058 1372
rect 4182 1368 4186 1372
rect 558 1358 562 1362
rect 910 1358 914 1362
rect 926 1358 930 1362
rect 1326 1358 1330 1362
rect 1334 1358 1338 1362
rect 1358 1358 1362 1362
rect 1374 1358 1378 1362
rect 1630 1358 1634 1362
rect 1758 1358 1762 1362
rect 1838 1358 1842 1362
rect 1886 1358 1890 1362
rect 1966 1358 1970 1362
rect 2014 1358 2018 1362
rect 2070 1358 2074 1362
rect 2318 1358 2322 1362
rect 2422 1358 2426 1362
rect 2590 1358 2594 1362
rect 2790 1358 2794 1362
rect 3214 1358 3218 1362
rect 3270 1358 3274 1362
rect 3542 1358 3546 1362
rect 3742 1358 3746 1362
rect 3782 1358 3786 1362
rect 4014 1358 4018 1362
rect 4118 1358 4122 1362
rect 4294 1358 4298 1362
rect 126 1348 130 1352
rect 710 1348 714 1352
rect 1062 1348 1066 1352
rect 1174 1348 1178 1352
rect 1270 1348 1274 1352
rect 1446 1348 1450 1352
rect 1486 1348 1490 1352
rect 1678 1348 1682 1352
rect 1734 1348 1738 1352
rect 1758 1348 1762 1352
rect 1774 1348 1778 1352
rect 1886 1348 1890 1352
rect 2334 1348 2338 1352
rect 2350 1348 2354 1352
rect 2550 1348 2554 1352
rect 3014 1348 3018 1352
rect 3278 1348 3282 1352
rect 3606 1348 3610 1352
rect 4126 1348 4130 1352
rect 4150 1348 4154 1352
rect 4182 1348 4186 1352
rect 4254 1348 4258 1352
rect 54 1338 58 1342
rect 246 1338 250 1342
rect 718 1338 722 1342
rect 886 1338 890 1342
rect 942 1338 946 1342
rect 1014 1338 1018 1342
rect 1134 1338 1138 1342
rect 1166 1338 1170 1342
rect 1230 1338 1234 1342
rect 1302 1338 1306 1342
rect 1374 1338 1378 1342
rect 1478 1338 1482 1342
rect 1582 1338 1586 1342
rect 1910 1338 1914 1342
rect 2294 1338 2298 1342
rect 3174 1338 3178 1342
rect 3246 1338 3250 1342
rect 3302 1338 3306 1342
rect 3350 1338 3354 1342
rect 3598 1338 3602 1342
rect 3646 1338 3650 1342
rect 3662 1338 3666 1342
rect 4310 1338 4314 1342
rect 758 1328 762 1332
rect 1414 1328 1418 1332
rect 2054 1328 2058 1332
rect 2606 1328 2610 1332
rect 2622 1328 2626 1332
rect 2638 1328 2642 1332
rect 2838 1328 2842 1332
rect 3286 1328 3290 1332
rect 3318 1328 3322 1332
rect 3326 1328 3330 1332
rect 3342 1328 3346 1332
rect 3542 1328 3546 1332
rect 3558 1328 3562 1332
rect 3782 1328 3786 1332
rect 4174 1328 4178 1332
rect 4254 1328 4258 1332
rect 662 1318 666 1322
rect 926 1318 930 1322
rect 1054 1318 1058 1322
rect 1486 1318 1490 1322
rect 1574 1318 1578 1322
rect 1606 1318 1610 1322
rect 1630 1318 1634 1322
rect 1694 1318 1698 1322
rect 1726 1318 1730 1322
rect 1742 1318 1746 1322
rect 1766 1318 1770 1322
rect 1798 1318 1802 1322
rect 1870 1318 1874 1322
rect 1878 1318 1882 1322
rect 2150 1318 2154 1322
rect 2406 1318 2410 1322
rect 3798 1318 3802 1322
rect 4230 1318 4234 1322
rect 694 1308 698 1312
rect 974 1308 978 1312
rect 1390 1308 1394 1312
rect 1486 1308 1490 1312
rect 1510 1308 1514 1312
rect 1566 1308 1570 1312
rect 1590 1308 1594 1312
rect 2086 1308 2090 1312
rect 2094 1308 2098 1312
rect 4382 1308 4386 1312
rect 898 1303 902 1307
rect 906 1303 909 1307
rect 909 1303 910 1307
rect 1930 1303 1934 1307
rect 1938 1303 1941 1307
rect 1941 1303 1942 1307
rect 2954 1303 2958 1307
rect 2962 1303 2965 1307
rect 2965 1303 2966 1307
rect 3978 1303 3982 1307
rect 3986 1303 3989 1307
rect 3989 1303 3990 1307
rect 6 1298 10 1302
rect 958 1298 962 1302
rect 1014 1298 1018 1302
rect 1382 1298 1386 1302
rect 2526 1298 2530 1302
rect 2534 1298 2538 1302
rect 3430 1298 3434 1302
rect 1070 1288 1074 1292
rect 1094 1288 1098 1292
rect 1110 1288 1114 1292
rect 1350 1288 1354 1292
rect 2038 1288 2042 1292
rect 2742 1288 2746 1292
rect 2974 1288 2978 1292
rect 3062 1288 3066 1292
rect 3222 1288 3226 1292
rect 3430 1288 3434 1292
rect 3750 1288 3754 1292
rect 4214 1288 4218 1292
rect 14 1278 18 1282
rect 142 1278 146 1282
rect 558 1278 562 1282
rect 726 1278 730 1282
rect 1086 1278 1090 1282
rect 1134 1278 1138 1282
rect 1206 1278 1210 1282
rect 1542 1278 1546 1282
rect 1822 1278 1826 1282
rect 2014 1278 2018 1282
rect 2062 1278 2066 1282
rect 2190 1278 2194 1282
rect 2222 1278 2226 1282
rect 2294 1278 2298 1282
rect 2406 1278 2410 1282
rect 2734 1278 2738 1282
rect 2798 1278 2802 1282
rect 3046 1278 3050 1282
rect 3166 1278 3170 1282
rect 3174 1278 3178 1282
rect 3398 1278 3402 1282
rect 3622 1278 3626 1282
rect 3678 1278 3682 1282
rect 3686 1278 3690 1282
rect 3878 1278 3882 1282
rect 4118 1278 4122 1282
rect 110 1268 114 1272
rect 534 1268 538 1272
rect 638 1268 642 1272
rect 646 1268 650 1272
rect 662 1268 666 1272
rect 974 1268 978 1272
rect 1070 1268 1074 1272
rect 1326 1268 1330 1272
rect 1334 1268 1338 1272
rect 1470 1268 1474 1272
rect 1598 1268 1602 1272
rect 1630 1268 1634 1272
rect 1758 1268 1762 1272
rect 2206 1268 2210 1272
rect 2286 1268 2290 1272
rect 2430 1268 2434 1272
rect 2606 1268 2610 1272
rect 2782 1268 2786 1272
rect 2902 1268 2906 1272
rect 3182 1268 3186 1272
rect 3222 1268 3226 1272
rect 3366 1268 3370 1272
rect 3430 1268 3434 1272
rect 3598 1268 3602 1272
rect 4222 1268 4226 1272
rect 4334 1268 4338 1272
rect 494 1258 498 1262
rect 526 1258 530 1262
rect 726 1258 730 1262
rect 822 1258 826 1262
rect 1134 1258 1138 1262
rect 1166 1258 1170 1262
rect 1182 1258 1186 1262
rect 1286 1258 1290 1262
rect 1334 1258 1338 1262
rect 1342 1258 1346 1262
rect 1422 1258 1426 1262
rect 1526 1258 1530 1262
rect 1534 1258 1538 1262
rect 1758 1258 1762 1262
rect 1766 1258 1770 1262
rect 1950 1258 1954 1262
rect 2502 1258 2506 1262
rect 2942 1258 2946 1262
rect 3150 1258 3154 1262
rect 3406 1258 3410 1262
rect 3758 1258 3762 1262
rect 3774 1258 3778 1262
rect 3910 1258 3914 1262
rect 4022 1258 4026 1262
rect 4158 1258 4162 1262
rect 14 1248 18 1252
rect 454 1248 458 1252
rect 574 1248 578 1252
rect 622 1248 626 1252
rect 678 1248 682 1252
rect 926 1248 930 1252
rect 950 1248 954 1252
rect 1494 1248 1498 1252
rect 1502 1248 1506 1252
rect 1630 1248 1634 1252
rect 1638 1248 1642 1252
rect 2590 1248 2594 1252
rect 3398 1248 3402 1252
rect 3646 1248 3650 1252
rect 3718 1248 3722 1252
rect 3870 1248 3874 1252
rect 4046 1248 4050 1252
rect 798 1238 802 1242
rect 846 1238 850 1242
rect 1158 1238 1162 1242
rect 1542 1238 1546 1242
rect 1654 1238 1658 1242
rect 1710 1238 1714 1242
rect 1750 1238 1754 1242
rect 2110 1238 2114 1242
rect 2686 1238 2690 1242
rect 3390 1238 3394 1242
rect 3582 1238 3586 1242
rect 4062 1238 4066 1242
rect 4238 1238 4242 1242
rect 686 1228 690 1232
rect 1566 1228 1570 1232
rect 1742 1228 1746 1232
rect 1750 1228 1754 1232
rect 1910 1228 1914 1232
rect 2142 1228 2146 1232
rect 3214 1228 3218 1232
rect 4142 1228 4146 1232
rect 926 1218 930 1222
rect 1110 1218 1114 1222
rect 1142 1218 1146 1222
rect 1606 1218 1610 1222
rect 1662 1218 1666 1222
rect 1862 1218 1866 1222
rect 2134 1218 2138 1222
rect 2622 1218 2626 1222
rect 2974 1218 2978 1222
rect 870 1208 874 1212
rect 1494 1208 1498 1212
rect 3238 1208 3242 1212
rect 3446 1208 3450 1212
rect 3526 1208 3530 1212
rect 394 1203 398 1207
rect 402 1203 405 1207
rect 405 1203 406 1207
rect 1418 1203 1422 1207
rect 1426 1203 1429 1207
rect 1429 1203 1430 1207
rect 2442 1203 2446 1207
rect 2450 1203 2453 1207
rect 2453 1203 2454 1207
rect 3474 1203 3478 1207
rect 3482 1203 3485 1207
rect 3485 1203 3486 1207
rect 118 1198 122 1202
rect 414 1198 418 1202
rect 566 1198 570 1202
rect 758 1198 762 1202
rect 982 1198 986 1202
rect 1550 1198 1554 1202
rect 1598 1198 1602 1202
rect 1974 1198 1978 1202
rect 3062 1198 3066 1202
rect 3302 1198 3306 1202
rect 3574 1198 3578 1202
rect 3606 1198 3610 1202
rect 3694 1198 3698 1202
rect 3862 1198 3866 1202
rect 3958 1198 3962 1202
rect 4286 1198 4290 1202
rect 6 1188 10 1192
rect 926 1188 930 1192
rect 1494 1188 1498 1192
rect 1894 1188 1898 1192
rect 2102 1188 2106 1192
rect 2590 1188 2594 1192
rect 3582 1188 3586 1192
rect 4198 1188 4202 1192
rect 14 1178 18 1182
rect 382 1178 386 1182
rect 702 1178 706 1182
rect 1430 1178 1434 1182
rect 1790 1178 1794 1182
rect 1854 1178 1858 1182
rect 1974 1178 1978 1182
rect 3078 1178 3082 1182
rect 3206 1178 3210 1182
rect 3462 1178 3466 1182
rect 3558 1178 3562 1182
rect 3566 1178 3570 1182
rect 3710 1178 3714 1182
rect 4054 1178 4058 1182
rect 94 1168 98 1172
rect 414 1168 418 1172
rect 1094 1168 1098 1172
rect 1358 1168 1362 1172
rect 1718 1168 1722 1172
rect 1758 1168 1762 1172
rect 1958 1168 1962 1172
rect 2262 1168 2266 1172
rect 2278 1168 2282 1172
rect 2854 1168 2858 1172
rect 2902 1168 2906 1172
rect 3166 1168 3170 1172
rect 3302 1168 3306 1172
rect 3750 1168 3754 1172
rect 3774 1168 3778 1172
rect 510 1158 514 1162
rect 766 1158 770 1162
rect 942 1158 946 1162
rect 1062 1158 1066 1162
rect 1102 1158 1106 1162
rect 1126 1158 1130 1162
rect 1358 1158 1362 1162
rect 1558 1158 1562 1162
rect 1662 1158 1666 1162
rect 1726 1158 1730 1162
rect 1918 1158 1922 1162
rect 2022 1158 2026 1162
rect 2214 1158 2218 1162
rect 2238 1158 2242 1162
rect 2574 1158 2578 1162
rect 2814 1158 2818 1162
rect 2822 1158 2826 1162
rect 3046 1158 3050 1162
rect 3054 1158 3058 1162
rect 3158 1158 3162 1162
rect 3694 1158 3698 1162
rect 3710 1158 3714 1162
rect 3998 1158 4002 1162
rect 4158 1158 4162 1162
rect 4222 1158 4226 1162
rect 4286 1158 4290 1162
rect 614 1148 618 1152
rect 678 1148 682 1152
rect 806 1148 810 1152
rect 926 1148 930 1152
rect 1070 1148 1074 1152
rect 1118 1148 1122 1152
rect 1142 1148 1146 1152
rect 1326 1148 1330 1152
rect 1334 1148 1338 1152
rect 1510 1148 1514 1152
rect 1694 1148 1698 1152
rect 1718 1148 1722 1152
rect 1998 1148 2002 1152
rect 2014 1148 2018 1152
rect 2126 1148 2130 1152
rect 2206 1148 2210 1152
rect 2222 1148 2226 1152
rect 2558 1148 2562 1152
rect 2878 1148 2882 1152
rect 3070 1148 3074 1152
rect 3102 1148 3106 1152
rect 3118 1148 3122 1152
rect 3142 1148 3146 1152
rect 3158 1148 3162 1152
rect 3254 1148 3258 1152
rect 3478 1148 3482 1152
rect 3502 1148 3506 1152
rect 3542 1148 3546 1152
rect 3630 1148 3634 1152
rect 3726 1148 3730 1152
rect 3782 1148 3786 1152
rect 4054 1148 4058 1152
rect 4294 1148 4298 1152
rect 374 1138 378 1142
rect 718 1138 722 1142
rect 982 1138 986 1142
rect 1230 1138 1234 1142
rect 1382 1138 1386 1142
rect 1470 1138 1474 1142
rect 1510 1138 1514 1142
rect 1862 1138 1866 1142
rect 3398 1138 3402 1142
rect 3614 1138 3618 1142
rect 3678 1138 3682 1142
rect 3758 1138 3762 1142
rect 270 1128 274 1132
rect 654 1128 658 1132
rect 782 1128 786 1132
rect 886 1128 890 1132
rect 1206 1128 1210 1132
rect 1230 1128 1234 1132
rect 1494 1128 1498 1132
rect 1534 1128 1538 1132
rect 1550 1128 1554 1132
rect 1814 1128 1818 1132
rect 1870 1128 1874 1132
rect 1958 1128 1962 1132
rect 2006 1128 2010 1132
rect 2198 1128 2202 1132
rect 2222 1128 2226 1132
rect 2398 1128 2402 1132
rect 2814 1128 2818 1132
rect 2990 1128 2994 1132
rect 3006 1128 3010 1132
rect 3086 1128 3090 1132
rect 3150 1128 3154 1132
rect 3198 1128 3202 1132
rect 3222 1128 3226 1132
rect 3502 1128 3506 1132
rect 3878 1128 3882 1132
rect 4302 1128 4306 1132
rect 294 1118 298 1122
rect 422 1118 426 1122
rect 798 1118 802 1122
rect 934 1118 938 1122
rect 1046 1118 1050 1122
rect 1206 1118 1210 1122
rect 1246 1118 1250 1122
rect 1350 1118 1354 1122
rect 1398 1118 1402 1122
rect 1622 1118 1626 1122
rect 1654 1118 1658 1122
rect 1678 1118 1682 1122
rect 1710 1118 1714 1122
rect 1918 1118 1922 1122
rect 2134 1118 2138 1122
rect 2254 1118 2258 1122
rect 2654 1118 2658 1122
rect 2742 1118 2746 1122
rect 2830 1118 2834 1122
rect 2998 1118 3002 1122
rect 3246 1118 3250 1122
rect 3390 1118 3394 1122
rect 3526 1118 3530 1122
rect 3694 1118 3698 1122
rect 4070 1118 4074 1122
rect 4086 1118 4090 1122
rect 4270 1118 4274 1122
rect 966 1108 970 1112
rect 1262 1108 1266 1112
rect 1374 1108 1378 1112
rect 1390 1108 1394 1112
rect 1822 1108 1826 1112
rect 2166 1108 2170 1112
rect 2198 1108 2202 1112
rect 2390 1108 2394 1112
rect 2422 1108 2426 1112
rect 2766 1108 2770 1112
rect 2862 1108 2866 1112
rect 2942 1108 2946 1112
rect 2982 1108 2986 1112
rect 3422 1108 3426 1112
rect 3718 1108 3722 1112
rect 4366 1108 4370 1112
rect 898 1103 902 1107
rect 906 1103 909 1107
rect 909 1103 910 1107
rect 1930 1103 1934 1107
rect 1938 1103 1941 1107
rect 1941 1103 1942 1107
rect 182 1098 186 1102
rect 678 1098 682 1102
rect 734 1098 738 1102
rect 862 1098 866 1102
rect 1470 1098 1474 1102
rect 1486 1098 1490 1102
rect 2954 1103 2958 1107
rect 2962 1103 2965 1107
rect 2965 1103 2966 1107
rect 3978 1103 3982 1107
rect 3986 1103 3989 1107
rect 3989 1103 3990 1107
rect 870 1088 874 1092
rect 1334 1088 1338 1092
rect 1526 1088 1530 1092
rect 1630 1088 1634 1092
rect 2398 1088 2402 1092
rect 2702 1088 2706 1092
rect 3542 1088 3546 1092
rect 3622 1088 3626 1092
rect 3710 1088 3714 1092
rect 4310 1088 4314 1092
rect 142 1078 146 1082
rect 438 1078 442 1082
rect 542 1078 546 1082
rect 766 1078 770 1082
rect 950 1078 954 1082
rect 1270 1078 1274 1082
rect 1566 1078 1570 1082
rect 1582 1078 1586 1082
rect 1766 1078 1770 1082
rect 1974 1078 1978 1082
rect 2030 1078 2034 1082
rect 2118 1078 2122 1082
rect 2318 1078 2322 1082
rect 2430 1078 2434 1082
rect 2534 1078 2538 1082
rect 2590 1078 2594 1082
rect 2774 1078 2778 1082
rect 2886 1078 2890 1082
rect 3094 1078 3098 1082
rect 3142 1078 3146 1082
rect 3206 1078 3210 1082
rect 3278 1078 3282 1082
rect 3286 1078 3290 1082
rect 3454 1078 3458 1082
rect 3574 1078 3578 1082
rect 3726 1078 3730 1082
rect 3742 1078 3746 1082
rect 3942 1078 3946 1082
rect 4190 1078 4194 1082
rect 4342 1078 4346 1082
rect 4390 1078 4394 1082
rect 158 1068 162 1072
rect 990 1068 994 1072
rect 998 1068 1002 1072
rect 1046 1068 1050 1072
rect 1070 1068 1074 1072
rect 1278 1068 1282 1072
rect 1302 1068 1306 1072
rect 414 1058 418 1062
rect 662 1058 666 1062
rect 750 1058 754 1062
rect 966 1058 970 1062
rect 982 1058 986 1062
rect 1078 1058 1082 1062
rect 1174 1058 1178 1062
rect 1406 1068 1410 1072
rect 1542 1068 1546 1072
rect 1774 1068 1778 1072
rect 1814 1068 1818 1072
rect 1854 1068 1858 1072
rect 1862 1068 1866 1072
rect 1950 1068 1954 1072
rect 2406 1068 2410 1072
rect 2550 1068 2554 1072
rect 2702 1068 2706 1072
rect 2934 1068 2938 1072
rect 2974 1068 2978 1072
rect 3110 1068 3114 1072
rect 3574 1068 3578 1072
rect 3742 1068 3746 1072
rect 3790 1068 3794 1072
rect 3958 1068 3962 1072
rect 4134 1068 4138 1072
rect 4198 1068 4202 1072
rect 4238 1068 4242 1072
rect 1462 1058 1466 1062
rect 1486 1058 1490 1062
rect 1566 1058 1570 1062
rect 1638 1058 1642 1062
rect 1646 1058 1650 1062
rect 1686 1058 1690 1062
rect 1726 1058 1730 1062
rect 2054 1058 2058 1062
rect 2942 1058 2946 1062
rect 3246 1058 3250 1062
rect 3470 1058 3474 1062
rect 3566 1058 3570 1062
rect 3598 1058 3602 1062
rect 3678 1058 3682 1062
rect 4062 1058 4066 1062
rect 4150 1058 4154 1062
rect 4166 1058 4170 1062
rect 4326 1058 4330 1062
rect 766 1048 770 1052
rect 862 1048 866 1052
rect 1150 1048 1154 1052
rect 1582 1048 1586 1052
rect 1590 1048 1594 1052
rect 1678 1048 1682 1052
rect 1806 1048 1810 1052
rect 1830 1048 1834 1052
rect 2094 1048 2098 1052
rect 2286 1048 2290 1052
rect 2318 1048 2322 1052
rect 2374 1048 2378 1052
rect 2478 1048 2482 1052
rect 2862 1048 2866 1052
rect 3358 1048 3362 1052
rect 4022 1048 4026 1052
rect 4158 1048 4162 1052
rect 4294 1048 4298 1052
rect 670 1038 674 1042
rect 1566 1038 1570 1042
rect 1870 1038 1874 1042
rect 3238 1038 3242 1042
rect 3598 1038 3602 1042
rect 3646 1038 3650 1042
rect 4246 1038 4250 1042
rect 4270 1038 4274 1042
rect 1142 1028 1146 1032
rect 1886 1028 1890 1032
rect 3574 1028 3578 1032
rect 3822 1028 3826 1032
rect 4102 1028 4106 1032
rect 4174 1028 4178 1032
rect 4222 1028 4226 1032
rect 1038 1018 1042 1022
rect 1062 1018 1066 1022
rect 1462 1018 1466 1022
rect 1574 1018 1578 1022
rect 1582 1018 1586 1022
rect 1942 1018 1946 1022
rect 2246 1018 2250 1022
rect 526 1008 530 1012
rect 686 1008 690 1012
rect 878 1008 882 1012
rect 1038 1008 1042 1012
rect 1166 1008 1170 1012
rect 1374 1008 1378 1012
rect 1878 1008 1882 1012
rect 1958 1008 1962 1012
rect 3022 1008 3026 1012
rect 3342 1008 3346 1012
rect 3622 1008 3626 1012
rect 3838 1008 3842 1012
rect 4070 1008 4074 1012
rect 394 1003 398 1007
rect 402 1003 405 1007
rect 405 1003 406 1007
rect 1418 1003 1422 1007
rect 1426 1003 1429 1007
rect 1429 1003 1430 1007
rect 2442 1003 2446 1007
rect 2450 1003 2453 1007
rect 2453 1003 2454 1007
rect 3474 1003 3478 1007
rect 3482 1003 3485 1007
rect 3485 1003 3486 1007
rect 1134 998 1138 1002
rect 1582 998 1586 1002
rect 1918 998 1922 1002
rect 3014 998 3018 1002
rect 294 988 298 992
rect 1654 988 1658 992
rect 1790 988 1794 992
rect 1990 988 1994 992
rect 2606 988 2610 992
rect 2638 988 2642 992
rect 3238 988 3242 992
rect 3718 998 3722 1002
rect 3630 988 3634 992
rect 4086 988 4090 992
rect 14 978 18 982
rect 1198 978 1202 982
rect 1318 978 1322 982
rect 2142 978 2146 982
rect 2358 978 2362 982
rect 2430 978 2434 982
rect 2742 978 2746 982
rect 2894 978 2898 982
rect 1166 968 1170 972
rect 1342 968 1346 972
rect 3454 968 3458 972
rect 3710 968 3714 972
rect 3718 968 3722 972
rect 4054 968 4058 972
rect 1102 958 1106 962
rect 1182 958 1186 962
rect 1206 958 1210 962
rect 1286 958 1290 962
rect 1326 958 1330 962
rect 1350 958 1354 962
rect 1438 958 1442 962
rect 1510 958 1514 962
rect 1558 958 1562 962
rect 1742 958 1746 962
rect 2022 958 2026 962
rect 2046 958 2050 962
rect 3318 958 3322 962
rect 3622 958 3626 962
rect 3958 958 3962 962
rect 4198 958 4202 962
rect 4214 958 4218 962
rect 4246 958 4250 962
rect 14 948 18 952
rect 542 948 546 952
rect 1054 948 1058 952
rect 1142 948 1146 952
rect 1158 948 1162 952
rect 1222 948 1226 952
rect 1230 948 1234 952
rect 1254 948 1258 952
rect 1270 948 1274 952
rect 1366 948 1370 952
rect 1758 948 1762 952
rect 1790 948 1794 952
rect 1870 948 1874 952
rect 2110 948 2114 952
rect 2502 948 2506 952
rect 2750 948 2754 952
rect 2774 948 2778 952
rect 3118 948 3122 952
rect 3134 948 3138 952
rect 590 938 594 942
rect 854 938 858 942
rect 1006 938 1010 942
rect 1046 938 1050 942
rect 1086 938 1090 942
rect 1134 938 1138 942
rect 1446 938 1450 942
rect 1494 938 1498 942
rect 1566 938 1570 942
rect 1822 938 1826 942
rect 1854 938 1858 942
rect 2062 938 2066 942
rect 2158 938 2162 942
rect 2526 938 2530 942
rect 2678 938 2682 942
rect 2886 938 2890 942
rect 3150 938 3154 942
rect 3390 948 3394 952
rect 3662 948 3666 952
rect 3766 948 3770 952
rect 4110 948 4114 952
rect 4182 948 4186 952
rect 3350 938 3354 942
rect 3414 938 3418 942
rect 3750 938 3754 942
rect 3774 938 3778 942
rect 3822 938 3826 942
rect 4118 938 4122 942
rect 4254 938 4258 942
rect 4262 938 4266 942
rect 4286 938 4290 942
rect 150 928 154 932
rect 374 928 378 932
rect 774 928 778 932
rect 1094 928 1098 932
rect 1606 928 1610 932
rect 1646 928 1650 932
rect 1702 928 1706 932
rect 1758 928 1762 932
rect 1854 928 1858 932
rect 1918 928 1922 932
rect 1942 928 1946 932
rect 2126 928 2130 932
rect 3294 928 3298 932
rect 3310 928 3314 932
rect 3422 928 3426 932
rect 846 918 850 922
rect 1038 918 1042 922
rect 1214 918 1218 922
rect 1342 918 1346 922
rect 1358 918 1362 922
rect 1558 918 1562 922
rect 1574 918 1578 922
rect 1638 918 1642 922
rect 1982 918 1986 922
rect 1990 918 1994 922
rect 2414 918 2418 922
rect 2918 918 2922 922
rect 3590 918 3594 922
rect 3910 918 3914 922
rect 4006 918 4010 922
rect 886 908 890 912
rect 942 908 946 912
rect 1126 908 1130 912
rect 1286 908 1290 912
rect 1502 908 1506 912
rect 1518 908 1522 912
rect 1886 908 1890 912
rect 1990 908 1994 912
rect 2390 908 2394 912
rect 2678 908 2682 912
rect 3086 908 3090 912
rect 3126 908 3130 912
rect 3998 908 4002 912
rect 4270 908 4274 912
rect 898 903 902 907
rect 906 903 909 907
rect 909 903 910 907
rect 1930 903 1934 907
rect 1938 903 1941 907
rect 1941 903 1942 907
rect 2954 903 2958 907
rect 2962 903 2965 907
rect 2965 903 2966 907
rect 3978 903 3982 907
rect 3986 903 3989 907
rect 3989 903 3990 907
rect 766 898 770 902
rect 854 898 858 902
rect 918 898 922 902
rect 1334 898 1338 902
rect 1390 898 1394 902
rect 1686 898 1690 902
rect 2046 898 2050 902
rect 2350 898 2354 902
rect 2942 898 2946 902
rect 3262 898 3266 902
rect 3526 898 3530 902
rect 774 888 778 892
rect 1110 888 1114 892
rect 1390 888 1394 892
rect 1462 888 1466 892
rect 1470 888 1474 892
rect 1718 888 1722 892
rect 3094 888 3098 892
rect 3126 888 3130 892
rect 3174 888 3178 892
rect 3542 888 3546 892
rect 3550 888 3554 892
rect 3718 888 3722 892
rect 3862 888 3866 892
rect 4190 888 4194 892
rect 422 878 426 882
rect 790 878 794 882
rect 814 878 818 882
rect 990 878 994 882
rect 1510 878 1514 882
rect 1622 878 1626 882
rect 1718 878 1722 882
rect 1798 878 1802 882
rect 1822 878 1826 882
rect 1846 878 1850 882
rect 1886 878 1890 882
rect 2086 878 2090 882
rect 2374 878 2378 882
rect 2590 878 2594 882
rect 2614 878 2618 882
rect 2662 878 2666 882
rect 158 868 162 872
rect 374 868 378 872
rect 766 868 770 872
rect 1014 868 1018 872
rect 1142 868 1146 872
rect 1678 868 1682 872
rect 1718 868 1722 872
rect 1734 868 1738 872
rect 1774 868 1778 872
rect 1974 868 1978 872
rect 2222 868 2226 872
rect 2310 868 2314 872
rect 2406 868 2410 872
rect 2766 868 2770 872
rect 2798 868 2802 872
rect 3662 878 3666 882
rect 3702 878 3706 882
rect 4150 878 4154 882
rect 4198 878 4202 882
rect 3182 868 3186 872
rect 3246 868 3250 872
rect 3846 868 3850 872
rect 4126 868 4130 872
rect 4206 868 4210 872
rect 4310 868 4314 872
rect 750 858 754 862
rect 822 858 826 862
rect 1038 858 1042 862
rect 1318 858 1322 862
rect 2406 858 2410 862
rect 2486 858 2490 862
rect 2630 858 2634 862
rect 2806 858 2810 862
rect 2894 858 2898 862
rect 3158 858 3162 862
rect 3238 858 3242 862
rect 3334 858 3338 862
rect 3406 858 3410 862
rect 3702 858 3706 862
rect 3710 858 3714 862
rect 3894 858 3898 862
rect 4190 858 4194 862
rect 4246 858 4250 862
rect 4286 858 4290 862
rect 518 848 522 852
rect 1382 848 1386 852
rect 1934 848 1938 852
rect 2622 848 2626 852
rect 2654 848 2658 852
rect 2886 848 2890 852
rect 2902 848 2906 852
rect 2926 848 2930 852
rect 2934 848 2938 852
rect 3022 848 3026 852
rect 3238 848 3242 852
rect 3926 848 3930 852
rect 4150 848 4154 852
rect 4286 848 4290 852
rect 4334 848 4338 852
rect 4366 848 4370 852
rect 702 838 706 842
rect 974 838 978 842
rect 1454 838 1458 842
rect 1590 838 1594 842
rect 1654 838 1658 842
rect 1670 838 1674 842
rect 1710 838 1714 842
rect 1790 838 1794 842
rect 2086 838 2090 842
rect 2974 838 2978 842
rect 3070 838 3074 842
rect 3190 838 3194 842
rect 3198 838 3202 842
rect 3286 838 3290 842
rect 3494 838 3498 842
rect 3894 838 3898 842
rect 1366 828 1370 832
rect 1782 828 1786 832
rect 1862 828 1866 832
rect 1902 828 1906 832
rect 2566 828 2570 832
rect 2902 828 2906 832
rect 3078 828 3082 832
rect 3166 828 3170 832
rect 3806 828 3810 832
rect 4150 828 4154 832
rect 1118 818 1122 822
rect 1398 818 1402 822
rect 2286 818 2290 822
rect 2598 818 2602 822
rect 2622 818 2626 822
rect 2822 818 2826 822
rect 2854 818 2858 822
rect 3838 818 3842 822
rect 4166 818 4170 822
rect 742 808 746 812
rect 1406 808 1410 812
rect 1638 808 1642 812
rect 1702 808 1706 812
rect 1806 808 1810 812
rect 2302 808 2306 812
rect 2662 808 2666 812
rect 3566 808 3570 812
rect 394 803 398 807
rect 402 803 405 807
rect 405 803 406 807
rect 1418 803 1422 807
rect 1426 803 1429 807
rect 1429 803 1430 807
rect 2442 803 2446 807
rect 2450 803 2453 807
rect 2453 803 2454 807
rect 3474 803 3478 807
rect 3482 803 3485 807
rect 3485 803 3486 807
rect 926 798 930 802
rect 1310 798 1314 802
rect 1494 798 1498 802
rect 1646 798 1650 802
rect 1862 798 1866 802
rect 2414 798 2418 802
rect 2670 798 2674 802
rect 2886 798 2890 802
rect 3206 798 3210 802
rect 3782 798 3786 802
rect 4054 798 4058 802
rect 4126 798 4130 802
rect 534 788 538 792
rect 734 788 738 792
rect 3294 788 3298 792
rect 4118 788 4122 792
rect 102 778 106 782
rect 430 778 434 782
rect 734 778 738 782
rect 806 778 810 782
rect 1598 778 1602 782
rect 2038 778 2042 782
rect 2294 778 2298 782
rect 2502 778 2506 782
rect 3118 778 3122 782
rect 3606 778 3610 782
rect 2270 768 2274 772
rect 2502 768 2506 772
rect 2854 768 2858 772
rect 3566 768 3570 772
rect 3622 768 3626 772
rect 3654 768 3658 772
rect 3726 768 3730 772
rect 4054 768 4058 772
rect 1118 758 1122 762
rect 1134 758 1138 762
rect 2030 758 2034 762
rect 2078 758 2082 762
rect 2190 758 2194 762
rect 2382 758 2386 762
rect 2910 758 2914 762
rect 2918 758 2922 762
rect 3462 758 3466 762
rect 3606 758 3610 762
rect 3614 758 3618 762
rect 3806 758 3810 762
rect 3822 758 3826 762
rect 3934 758 3938 762
rect 4062 758 4066 762
rect 4110 758 4114 762
rect 4198 758 4202 762
rect 726 748 730 752
rect 982 748 986 752
rect 1126 748 1130 752
rect 1190 748 1194 752
rect 1430 748 1434 752
rect 1454 748 1458 752
rect 1694 748 1698 752
rect 1702 748 1706 752
rect 1734 748 1738 752
rect 1742 748 1746 752
rect 1966 748 1970 752
rect 2014 748 2018 752
rect 2046 748 2050 752
rect 2350 748 2354 752
rect 2526 748 2530 752
rect 2566 748 2570 752
rect 2638 748 2642 752
rect 2678 748 2682 752
rect 3382 748 3386 752
rect 3646 748 3650 752
rect 3718 748 3722 752
rect 3846 748 3850 752
rect 4062 748 4066 752
rect 4118 748 4122 752
rect 4270 748 4274 752
rect 4382 748 4386 752
rect 158 738 162 742
rect 574 738 578 742
rect 734 738 738 742
rect 918 738 922 742
rect 1070 738 1074 742
rect 1334 738 1338 742
rect 1366 738 1370 742
rect 1462 738 1466 742
rect 1494 738 1498 742
rect 1718 738 1722 742
rect 1798 738 1802 742
rect 2174 738 2178 742
rect 2230 738 2234 742
rect 2302 738 2306 742
rect 2358 738 2362 742
rect 2398 738 2402 742
rect 2510 738 2514 742
rect 2598 738 2602 742
rect 3302 738 3306 742
rect 3502 738 3506 742
rect 3638 738 3642 742
rect 3830 738 3834 742
rect 3910 738 3914 742
rect 4246 738 4250 742
rect 726 728 730 732
rect 854 728 858 732
rect 1438 728 1442 732
rect 1838 728 1842 732
rect 1950 728 1954 732
rect 1438 718 1442 722
rect 1470 718 1474 722
rect 1614 718 1618 722
rect 1646 718 1650 722
rect 1654 718 1658 722
rect 1806 718 1810 722
rect 1814 718 1818 722
rect 1830 718 1834 722
rect 2526 728 2530 732
rect 2550 728 2554 732
rect 2750 728 2754 732
rect 2758 728 2762 732
rect 3110 728 3114 732
rect 3542 728 3546 732
rect 3710 728 3714 732
rect 3862 728 3866 732
rect 2158 718 2162 722
rect 2190 718 2194 722
rect 2518 718 2522 722
rect 2726 718 2730 722
rect 3174 718 3178 722
rect 3518 718 3522 722
rect 702 708 706 712
rect 1422 708 1426 712
rect 1614 708 1618 712
rect 1662 708 1666 712
rect 2110 708 2114 712
rect 2694 708 2698 712
rect 2878 708 2882 712
rect 2974 708 2978 712
rect 3246 708 3250 712
rect 4230 708 4234 712
rect 898 703 902 707
rect 906 703 909 707
rect 909 703 910 707
rect 1930 703 1934 707
rect 1938 703 1941 707
rect 1941 703 1942 707
rect 2954 703 2958 707
rect 2962 703 2965 707
rect 2965 703 2966 707
rect 3978 703 3982 707
rect 3986 703 3989 707
rect 3989 703 3990 707
rect 710 698 714 702
rect 918 698 922 702
rect 1078 698 1082 702
rect 1102 698 1106 702
rect 1326 698 1330 702
rect 1558 698 1562 702
rect 1694 698 1698 702
rect 2190 698 2194 702
rect 2310 698 2314 702
rect 2990 698 2994 702
rect 3358 698 3362 702
rect 3414 698 3418 702
rect 3438 698 3442 702
rect 3870 698 3874 702
rect 3902 698 3906 702
rect 254 688 258 692
rect 646 688 650 692
rect 518 678 522 682
rect 582 678 586 682
rect 1094 688 1098 692
rect 1782 688 1786 692
rect 1846 688 1850 692
rect 2318 688 2322 692
rect 2622 688 2626 692
rect 2894 688 2898 692
rect 3262 688 3266 692
rect 3366 688 3370 692
rect 3414 688 3418 692
rect 3630 688 3634 692
rect 3686 688 3690 692
rect 1446 678 1450 682
rect 1598 678 1602 682
rect 1870 678 1874 682
rect 1878 678 1882 682
rect 1926 678 1930 682
rect 2622 678 2626 682
rect 2798 678 2802 682
rect 3878 678 3882 682
rect 134 668 138 672
rect 382 668 386 672
rect 694 668 698 672
rect 1030 668 1034 672
rect 1230 668 1234 672
rect 1462 668 1466 672
rect 1486 668 1490 672
rect 1518 668 1522 672
rect 1894 668 1898 672
rect 2046 668 2050 672
rect 2110 668 2114 672
rect 2310 668 2314 672
rect 2918 668 2922 672
rect 3070 668 3074 672
rect 3374 668 3378 672
rect 3702 668 3706 672
rect 4022 668 4026 672
rect 4310 668 4314 672
rect 4358 668 4362 672
rect 846 658 850 662
rect 1398 658 1402 662
rect 1510 658 1514 662
rect 1606 658 1610 662
rect 1622 658 1626 662
rect 1670 658 1674 662
rect 1958 658 1962 662
rect 2582 658 2586 662
rect 2718 658 2722 662
rect 2990 658 2994 662
rect 3006 658 3010 662
rect 3358 658 3362 662
rect 3398 658 3402 662
rect 3454 658 3458 662
rect 3782 658 3786 662
rect 4214 658 4218 662
rect 4278 658 4282 662
rect 1222 648 1226 652
rect 1254 648 1258 652
rect 1318 648 1322 652
rect 1478 648 1482 652
rect 1566 648 1570 652
rect 1758 648 1762 652
rect 1766 648 1770 652
rect 1878 648 1882 652
rect 2990 648 2994 652
rect 3262 648 3266 652
rect 3286 648 3290 652
rect 3614 648 3618 652
rect 3774 648 3778 652
rect 3902 648 3906 652
rect 4078 648 4082 652
rect 4302 648 4306 652
rect 1022 638 1026 642
rect 1078 638 1082 642
rect 1710 638 1714 642
rect 2206 638 2210 642
rect 2238 638 2242 642
rect 2414 638 2418 642
rect 2630 638 2634 642
rect 3502 638 3506 642
rect 4046 638 4050 642
rect 4062 638 4066 642
rect 110 628 114 632
rect 1206 628 1210 632
rect 1574 628 1578 632
rect 2902 628 2906 632
rect 2998 628 3002 632
rect 3078 628 3082 632
rect 3350 628 3354 632
rect 270 618 274 622
rect 286 618 290 622
rect 1926 618 1930 622
rect 3598 618 3602 622
rect 94 608 98 612
rect 1366 608 1370 612
rect 2238 608 2242 612
rect 2422 608 2426 612
rect 2654 608 2658 612
rect 3238 608 3242 612
rect 3406 608 3410 612
rect 3598 608 3602 612
rect 3958 608 3962 612
rect 4366 608 4370 612
rect 394 603 398 607
rect 402 603 405 607
rect 405 603 406 607
rect 1418 603 1422 607
rect 1426 603 1429 607
rect 1429 603 1430 607
rect 2442 603 2446 607
rect 2450 603 2453 607
rect 2453 603 2454 607
rect 3474 603 3478 607
rect 3482 603 3485 607
rect 3485 603 3486 607
rect 1118 598 1122 602
rect 1126 598 1130 602
rect 2494 598 2498 602
rect 2774 598 2778 602
rect 3566 598 3570 602
rect 1078 588 1082 592
rect 1734 588 1738 592
rect 1974 588 1978 592
rect 2222 588 2226 592
rect 2422 588 2426 592
rect 2590 588 2594 592
rect 2894 588 2898 592
rect 3158 588 3162 592
rect 3214 588 3218 592
rect 3302 588 3306 592
rect 3614 588 3618 592
rect 3726 588 3730 592
rect 3798 588 3802 592
rect 438 578 442 582
rect 1438 578 1442 582
rect 2542 578 2546 582
rect 3566 578 3570 582
rect 3790 578 3794 582
rect 414 568 418 572
rect 1406 568 1410 572
rect 1462 568 1466 572
rect 1638 568 1642 572
rect 1862 568 1866 572
rect 1974 568 1978 572
rect 2022 568 2026 572
rect 2102 568 2106 572
rect 2174 568 2178 572
rect 2206 568 2210 572
rect 2654 568 2658 572
rect 3326 568 3330 572
rect 3518 568 3522 572
rect 3894 568 3898 572
rect 4086 568 4090 572
rect 4190 568 4194 572
rect 4230 568 4234 572
rect 4342 568 4346 572
rect 446 558 450 562
rect 1094 558 1098 562
rect 1270 558 1274 562
rect 2606 558 2610 562
rect 2686 558 2690 562
rect 2710 558 2714 562
rect 2830 558 2834 562
rect 3118 558 3122 562
rect 3174 558 3178 562
rect 3342 558 3346 562
rect 3902 558 3906 562
rect 4078 558 4082 562
rect 4110 558 4114 562
rect 4142 558 4146 562
rect 4174 558 4178 562
rect 4334 558 4338 562
rect 182 548 186 552
rect 958 548 962 552
rect 974 548 978 552
rect 1286 548 1290 552
rect 1422 548 1426 552
rect 1662 548 1666 552
rect 1806 548 1810 552
rect 2582 548 2586 552
rect 3462 548 3466 552
rect 3518 548 3522 552
rect 3934 548 3938 552
rect 4022 548 4026 552
rect 4262 548 4266 552
rect 4270 548 4274 552
rect 1102 538 1106 542
rect 1110 538 1114 542
rect 1286 538 1290 542
rect 1446 538 1450 542
rect 1478 538 1482 542
rect 1518 538 1522 542
rect 1982 538 1986 542
rect 2158 538 2162 542
rect 3206 538 3210 542
rect 3774 538 3778 542
rect 3870 538 3874 542
rect 4286 538 4290 542
rect 150 528 154 532
rect 566 528 570 532
rect 1214 528 1218 532
rect 1238 528 1242 532
rect 1558 528 1562 532
rect 1678 528 1682 532
rect 1758 528 1762 532
rect 1782 528 1786 532
rect 2006 528 2010 532
rect 2870 528 2874 532
rect 3254 528 3258 532
rect 3422 528 3426 532
rect 3918 528 3922 532
rect 4270 528 4274 532
rect 718 518 722 522
rect 886 518 890 522
rect 1246 518 1250 522
rect 1254 518 1258 522
rect 1390 518 1394 522
rect 1614 518 1618 522
rect 2022 518 2026 522
rect 2678 518 2682 522
rect 2774 518 2778 522
rect 3198 518 3202 522
rect 918 508 922 512
rect 998 508 1002 512
rect 1134 508 1138 512
rect 1774 508 1778 512
rect 2014 508 2018 512
rect 2654 508 2658 512
rect 2670 508 2674 512
rect 3294 508 3298 512
rect 898 503 902 507
rect 906 503 909 507
rect 909 503 910 507
rect 1930 503 1934 507
rect 1938 503 1941 507
rect 1941 503 1942 507
rect 2954 503 2958 507
rect 2962 503 2965 507
rect 2965 503 2966 507
rect 3978 503 3982 507
rect 3986 503 3989 507
rect 3989 503 3990 507
rect 1742 498 1746 502
rect 2550 498 2554 502
rect 2758 498 2762 502
rect 4054 498 4058 502
rect 1238 488 1242 492
rect 1582 488 1586 492
rect 1702 488 1706 492
rect 1998 488 2002 492
rect 2262 488 2266 492
rect 2350 488 2354 492
rect 2478 488 2482 492
rect 2958 488 2962 492
rect 3166 488 3170 492
rect 3350 488 3354 492
rect 3694 488 3698 492
rect 3814 488 3818 492
rect 142 478 146 482
rect 534 478 538 482
rect 1222 478 1226 482
rect 1262 478 1266 482
rect 1270 478 1274 482
rect 1302 478 1306 482
rect 1486 478 1490 482
rect 1606 478 1610 482
rect 2006 478 2010 482
rect 2054 478 2058 482
rect 2150 478 2154 482
rect 3158 478 3162 482
rect 3174 478 3178 482
rect 3550 478 3554 482
rect 3598 478 3602 482
rect 4006 478 4010 482
rect 1150 468 1154 472
rect 1446 468 1450 472
rect 1454 468 1458 472
rect 1494 468 1498 472
rect 1574 468 1578 472
rect 1998 468 2002 472
rect 2374 468 2378 472
rect 2462 468 2466 472
rect 2974 468 2978 472
rect 3118 468 3122 472
rect 3182 468 3186 472
rect 3310 468 3314 472
rect 3598 468 3602 472
rect 4006 468 4010 472
rect 710 458 714 462
rect 1366 458 1370 462
rect 1518 458 1522 462
rect 1526 458 1530 462
rect 1534 458 1538 462
rect 2342 458 2346 462
rect 2358 458 2362 462
rect 2774 458 2778 462
rect 3054 458 3058 462
rect 3094 458 3098 462
rect 3166 458 3170 462
rect 3230 458 3234 462
rect 3726 458 3730 462
rect 3822 458 3826 462
rect 4086 458 4090 462
rect 4190 458 4194 462
rect 1134 448 1138 452
rect 1838 448 1842 452
rect 2030 448 2034 452
rect 2110 448 2114 452
rect 2310 448 2314 452
rect 2510 448 2514 452
rect 2526 448 2530 452
rect 2558 448 2562 452
rect 2926 448 2930 452
rect 3022 448 3026 452
rect 4078 448 4082 452
rect 4118 448 4122 452
rect 4334 448 4338 452
rect 414 438 418 442
rect 558 438 562 442
rect 790 438 794 442
rect 1550 438 1554 442
rect 2334 438 2338 442
rect 2342 438 2346 442
rect 3094 438 3098 442
rect 3678 438 3682 442
rect 4214 438 4218 442
rect 4238 438 4242 442
rect 1118 428 1122 432
rect 2246 428 2250 432
rect 4102 428 4106 432
rect 4150 428 4154 432
rect 4302 428 4306 432
rect 118 418 122 422
rect 678 418 682 422
rect 854 418 858 422
rect 1174 418 1178 422
rect 1366 418 1370 422
rect 2102 418 2106 422
rect 2134 418 2138 422
rect 2486 418 2490 422
rect 3838 418 3842 422
rect 118 408 122 412
rect 918 408 922 412
rect 1230 408 1234 412
rect 1382 408 1386 412
rect 1878 408 1882 412
rect 2422 408 2426 412
rect 2566 408 2570 412
rect 3214 408 3218 412
rect 3494 408 3498 412
rect 394 403 398 407
rect 402 403 405 407
rect 405 403 406 407
rect 1418 403 1422 407
rect 1426 403 1429 407
rect 1429 403 1430 407
rect 2442 403 2446 407
rect 2450 403 2453 407
rect 2453 403 2454 407
rect 3474 403 3478 407
rect 3482 403 3485 407
rect 3485 403 3486 407
rect 766 398 770 402
rect 1646 398 1650 402
rect 1702 398 1706 402
rect 2238 398 2242 402
rect 2654 398 2658 402
rect 3742 398 3746 402
rect 3894 398 3898 402
rect 4174 398 4178 402
rect 550 388 554 392
rect 782 388 786 392
rect 790 388 794 392
rect 1230 388 1234 392
rect 2030 388 2034 392
rect 2126 388 2130 392
rect 2486 388 2490 392
rect 2646 388 2650 392
rect 2766 388 2770 392
rect 3062 388 3066 392
rect 3278 388 3282 392
rect 3326 388 3330 392
rect 4262 388 4266 392
rect 110 378 114 382
rect 982 378 986 382
rect 1798 378 1802 382
rect 1806 378 1810 382
rect 1918 378 1922 382
rect 1998 378 2002 382
rect 2102 378 2106 382
rect 2830 378 2834 382
rect 3710 378 3714 382
rect 3854 378 3858 382
rect 3886 378 3890 382
rect 4358 378 4362 382
rect 1310 368 1314 372
rect 1494 368 1498 372
rect 1894 368 1898 372
rect 2006 368 2010 372
rect 2302 368 2306 372
rect 2406 368 2410 372
rect 2526 368 2530 372
rect 3798 368 3802 372
rect 3934 368 3938 372
rect 182 358 186 362
rect 1182 358 1186 362
rect 1542 358 1546 362
rect 1590 358 1594 362
rect 2054 358 2058 362
rect 2230 358 2234 362
rect 2894 358 2898 362
rect 2990 358 2994 362
rect 3230 358 3234 362
rect 3494 358 3498 362
rect 3694 358 3698 362
rect 4062 358 4066 362
rect 4206 358 4210 362
rect 4238 358 4242 362
rect 4286 358 4290 362
rect 382 348 386 352
rect 710 348 714 352
rect 974 348 978 352
rect 1278 348 1282 352
rect 1894 348 1898 352
rect 2262 348 2266 352
rect 2390 348 2394 352
rect 2518 348 2522 352
rect 2574 348 2578 352
rect 3054 348 3058 352
rect 3262 348 3266 352
rect 3382 348 3386 352
rect 3462 348 3466 352
rect 3614 348 3618 352
rect 3822 348 3826 352
rect 3926 348 3930 352
rect 4030 348 4034 352
rect 4278 348 4282 352
rect 206 338 210 342
rect 886 338 890 342
rect 1070 338 1074 342
rect 1238 338 1242 342
rect 1550 338 1554 342
rect 1726 338 1730 342
rect 1886 338 1890 342
rect 1942 338 1946 342
rect 2046 338 2050 342
rect 2246 338 2250 342
rect 2862 338 2866 342
rect 3246 338 3250 342
rect 3718 338 3722 342
rect 3750 338 3754 342
rect 3910 338 3914 342
rect 3958 338 3962 342
rect 1150 328 1154 332
rect 1206 328 1210 332
rect 1214 328 1218 332
rect 1294 328 1298 332
rect 2086 328 2090 332
rect 2118 328 2122 332
rect 3518 328 3522 332
rect 3966 328 3970 332
rect 3974 328 3978 332
rect 358 318 362 322
rect 718 318 722 322
rect 1246 318 1250 322
rect 1334 318 1338 322
rect 1782 318 1786 322
rect 1830 318 1834 322
rect 1838 318 1842 322
rect 2398 318 2402 322
rect 3686 318 3690 322
rect 782 308 786 312
rect 918 308 922 312
rect 1758 308 1762 312
rect 2942 308 2946 312
rect 3958 308 3962 312
rect 4070 308 4074 312
rect 4374 308 4378 312
rect 898 303 902 307
rect 906 303 909 307
rect 909 303 910 307
rect 1930 303 1934 307
rect 1938 303 1941 307
rect 1941 303 1942 307
rect 2954 303 2958 307
rect 2962 303 2965 307
rect 2965 303 2966 307
rect 3978 303 3982 307
rect 3986 303 3989 307
rect 3989 303 3990 307
rect 1006 298 1010 302
rect 1262 298 1266 302
rect 1470 298 1474 302
rect 1670 298 1674 302
rect 1678 298 1682 302
rect 2118 298 2122 302
rect 2838 298 2842 302
rect 2926 298 2930 302
rect 3966 298 3970 302
rect 382 288 386 292
rect 542 288 546 292
rect 950 288 954 292
rect 1838 288 1842 292
rect 1990 288 1994 292
rect 2262 288 2266 292
rect 2358 288 2362 292
rect 2558 288 2562 292
rect 2566 288 2570 292
rect 2814 288 2818 292
rect 3054 288 3058 292
rect 3134 288 3138 292
rect 3406 288 3410 292
rect 3454 288 3458 292
rect 3742 288 3746 292
rect 4254 288 4258 292
rect 518 278 522 282
rect 1110 278 1114 282
rect 1590 278 1594 282
rect 1606 278 1610 282
rect 2270 278 2274 282
rect 2702 278 2706 282
rect 3102 278 3106 282
rect 3174 278 3178 282
rect 3590 278 3594 282
rect 3654 278 3658 282
rect 3926 278 3930 282
rect 110 268 114 272
rect 478 268 482 272
rect 534 268 538 272
rect 630 268 634 272
rect 1062 268 1066 272
rect 1230 268 1234 272
rect 1446 268 1450 272
rect 1486 268 1490 272
rect 1518 268 1522 272
rect 1982 268 1986 272
rect 2134 268 2138 272
rect 2374 268 2378 272
rect 2806 268 2810 272
rect 2934 268 2938 272
rect 3926 268 3930 272
rect 4086 268 4090 272
rect 4174 268 4178 272
rect 422 258 426 262
rect 1246 258 1250 262
rect 1350 258 1354 262
rect 1494 258 1498 262
rect 3174 258 3178 262
rect 3590 258 3594 262
rect 3894 258 3898 262
rect 4222 258 4226 262
rect 4302 258 4306 262
rect 838 248 842 252
rect 1230 248 1234 252
rect 1598 248 1602 252
rect 1718 248 1722 252
rect 2286 248 2290 252
rect 2334 248 2338 252
rect 2358 248 2362 252
rect 2414 248 2418 252
rect 2862 248 2866 252
rect 3102 248 3106 252
rect 3470 248 3474 252
rect 3638 248 3642 252
rect 4014 248 4018 252
rect 1326 238 1330 242
rect 2510 238 2514 242
rect 3054 238 3058 242
rect 1478 228 1482 232
rect 2094 228 2098 232
rect 2462 228 2466 232
rect 2550 228 2554 232
rect 3142 228 3146 232
rect 3822 228 3826 232
rect 3894 228 3898 232
rect 4118 228 4122 232
rect 4262 228 4266 232
rect 678 218 682 222
rect 1118 218 1122 222
rect 1390 218 1394 222
rect 1526 218 1530 222
rect 2038 218 2042 222
rect 3518 218 3522 222
rect 3710 218 3714 222
rect 3718 218 3722 222
rect 3886 218 3890 222
rect 1438 208 1442 212
rect 2118 208 2122 212
rect 2462 208 2466 212
rect 2942 208 2946 212
rect 2974 208 2978 212
rect 3710 208 3714 212
rect 3726 208 3730 212
rect 3734 208 3738 212
rect 3830 208 3834 212
rect 4198 208 4202 212
rect 394 203 398 207
rect 402 203 405 207
rect 405 203 406 207
rect 1418 203 1422 207
rect 1426 203 1429 207
rect 1429 203 1430 207
rect 2442 203 2446 207
rect 2450 203 2453 207
rect 2453 203 2454 207
rect 3474 203 3478 207
rect 3482 203 3485 207
rect 3485 203 3486 207
rect 1214 198 1218 202
rect 3358 198 3362 202
rect 3902 198 3906 202
rect 1198 188 1202 192
rect 1302 188 1306 192
rect 1398 188 1402 192
rect 2262 188 2266 192
rect 3246 188 3250 192
rect 3454 188 3458 192
rect 3918 188 3922 192
rect 374 178 378 182
rect 1262 178 1266 182
rect 2006 178 2010 182
rect 2326 178 2330 182
rect 2526 178 2530 182
rect 2654 178 2658 182
rect 3118 178 3122 182
rect 4294 178 4298 182
rect 4342 178 4346 182
rect 974 168 978 172
rect 3422 168 3426 172
rect 3462 168 3466 172
rect 4070 168 4074 172
rect 358 158 362 162
rect 990 158 994 162
rect 1182 158 1186 162
rect 1246 158 1250 162
rect 1270 158 1274 162
rect 1566 158 1570 162
rect 1934 158 1938 162
rect 2054 158 2058 162
rect 2358 158 2362 162
rect 3358 158 3362 162
rect 4302 158 4306 162
rect 4358 158 4362 162
rect 222 148 226 152
rect 974 148 978 152
rect 1374 148 1378 152
rect 1406 148 1410 152
rect 1550 148 1554 152
rect 1614 148 1618 152
rect 2038 148 2042 152
rect 2694 148 2698 152
rect 2710 148 2714 152
rect 2718 148 2722 152
rect 3814 148 3818 152
rect 4142 148 4146 152
rect 4294 148 4298 152
rect 254 138 258 142
rect 494 138 498 142
rect 694 138 698 142
rect 1030 138 1034 142
rect 1110 138 1114 142
rect 1158 138 1162 142
rect 1254 138 1258 142
rect 1318 138 1322 142
rect 1646 138 1650 142
rect 1718 138 1722 142
rect 2070 138 2074 142
rect 2078 138 2082 142
rect 2118 138 2122 142
rect 2222 138 2226 142
rect 2430 138 2434 142
rect 2494 138 2498 142
rect 3838 138 3842 142
rect 3862 138 3866 142
rect 3926 138 3930 142
rect 4318 138 4322 142
rect 1038 128 1042 132
rect 1094 128 1098 132
rect 1414 128 1418 132
rect 1710 128 1714 132
rect 1726 128 1730 132
rect 2014 128 2018 132
rect 2046 128 2050 132
rect 2350 128 2354 132
rect 2542 128 2546 132
rect 2558 128 2562 132
rect 3654 128 3658 132
rect 3742 128 3746 132
rect 3798 128 3802 132
rect 4302 128 4306 132
rect 4318 128 4322 132
rect 1334 118 1338 122
rect 1342 118 1346 122
rect 1654 118 1658 122
rect 2214 118 2218 122
rect 3182 118 3186 122
rect 3806 118 3810 122
rect 4102 118 4106 122
rect 286 108 290 112
rect 1286 108 1290 112
rect 1806 108 1810 112
rect 2334 108 2338 112
rect 2358 108 2362 112
rect 4038 108 4042 112
rect 4094 108 4098 112
rect 898 103 902 107
rect 906 103 909 107
rect 909 103 910 107
rect 1930 103 1934 107
rect 1938 103 1941 107
rect 1941 103 1942 107
rect 574 98 578 102
rect 774 98 778 102
rect 1382 98 1386 102
rect 1518 98 1522 102
rect 1734 98 1738 102
rect 2006 98 2010 102
rect 2954 103 2958 107
rect 2962 103 2965 107
rect 2965 103 2966 107
rect 3978 103 3982 107
rect 3986 103 3989 107
rect 3989 103 3990 107
rect 2806 98 2810 102
rect 3374 98 3378 102
rect 3798 98 3802 102
rect 4158 98 4162 102
rect 550 88 554 92
rect 1022 88 1026 92
rect 1358 88 1362 92
rect 1398 88 1402 92
rect 1670 88 1674 92
rect 2086 88 2090 92
rect 2606 88 2610 92
rect 3350 88 3354 92
rect 3566 88 3570 92
rect 3590 88 3594 92
rect 3726 88 3730 92
rect 4142 88 4146 92
rect 4150 88 4154 92
rect 4206 88 4210 92
rect 358 78 362 82
rect 478 78 482 82
rect 1038 78 1042 82
rect 1246 78 1250 82
rect 1510 78 1514 82
rect 2046 78 2050 82
rect 2126 78 2130 82
rect 2302 78 2306 82
rect 2670 78 2674 82
rect 2974 78 2978 82
rect 3078 78 3082 82
rect 3806 78 3810 82
rect 3902 78 3906 82
rect 4382 78 4386 82
rect 158 68 162 72
rect 254 68 258 72
rect 550 68 554 72
rect 1030 68 1034 72
rect 1102 68 1106 72
rect 1326 68 1330 72
rect 1374 68 1378 72
rect 1502 68 1506 72
rect 1734 68 1738 72
rect 2054 68 2058 72
rect 2238 68 2242 72
rect 2974 68 2978 72
rect 3678 68 3682 72
rect 3726 68 3730 72
rect 4182 68 4186 72
rect 4326 68 4330 72
rect 3174 58 3178 62
rect 3998 58 4002 62
rect 4134 58 4138 62
rect 4310 58 4314 62
rect 1022 48 1026 52
rect 1230 48 1234 52
rect 1598 48 1602 52
rect 2006 48 2010 52
rect 3374 48 3378 52
rect 4174 48 4178 52
rect 4166 38 4170 42
rect 1326 28 1330 32
rect 2286 28 2290 32
rect 542 18 546 22
rect 558 18 562 22
rect 1414 18 1418 22
rect 2094 18 2098 22
rect 350 8 354 12
rect 566 8 570 12
rect 638 8 642 12
rect 766 8 770 12
rect 1014 8 1018 12
rect 1190 8 1194 12
rect 1366 8 1370 12
rect 2158 8 2162 12
rect 2174 8 2178 12
rect 2502 8 2506 12
rect 2630 8 2634 12
rect 2742 8 2746 12
rect 394 3 398 7
rect 402 3 405 7
rect 405 3 406 7
rect 1418 3 1422 7
rect 1426 3 1429 7
rect 1429 3 1430 7
rect 2442 3 2446 7
rect 2450 3 2453 7
rect 2453 3 2454 7
rect 3474 3 3478 7
rect 3482 3 3485 7
rect 3485 3 3486 7
<< metal4 >>
rect 896 3103 898 3107
rect 902 3103 905 3107
rect 910 3103 912 3107
rect 1928 3103 1930 3107
rect 1934 3103 1937 3107
rect 1942 3103 1944 3107
rect 2952 3103 2954 3107
rect 2958 3103 2961 3107
rect 2966 3103 2968 3107
rect 3976 3103 3978 3107
rect 3982 3103 3985 3107
rect 3990 3103 3992 3107
rect 1134 3098 1142 3101
rect 1694 3098 1702 3101
rect 1898 3098 1905 3101
rect 630 3072 633 3078
rect 218 3068 222 3071
rect 314 3058 318 3061
rect 102 2872 105 3018
rect 392 3003 394 3007
rect 398 3003 401 3007
rect 406 3003 408 3007
rect 30 2742 33 2788
rect 38 2452 41 2588
rect 86 2482 89 2758
rect 94 2602 97 2708
rect 86 2332 89 2478
rect 26 2148 30 2151
rect 6 1952 9 1998
rect 70 1951 73 1958
rect 66 1948 73 1951
rect 10 1788 14 1791
rect 6 1622 9 1648
rect 6 1492 9 1508
rect 14 1492 17 1548
rect 102 1542 105 2868
rect 214 2642 217 2758
rect 114 2558 118 2561
rect 166 2082 169 2278
rect 174 2132 177 2338
rect 182 2142 185 2168
rect 194 2148 198 2151
rect 206 1952 209 2118
rect 162 1938 166 1941
rect 162 1738 166 1741
rect 158 1672 161 1678
rect 166 1662 169 1678
rect 174 1552 177 1948
rect 186 1938 190 1941
rect 334 1932 337 2498
rect 382 2332 385 2898
rect 550 2862 553 3068
rect 706 3058 710 3061
rect 726 3038 734 3041
rect 392 2803 394 2807
rect 398 2803 401 2807
rect 406 2803 408 2807
rect 526 2742 529 2808
rect 534 2792 537 2838
rect 392 2603 394 2607
rect 398 2603 401 2607
rect 406 2603 408 2607
rect 392 2403 394 2407
rect 398 2403 401 2407
rect 406 2403 408 2407
rect 366 2042 369 2318
rect 392 2203 394 2207
rect 398 2203 401 2207
rect 406 2203 408 2207
rect 422 2202 425 2728
rect 534 2662 537 2748
rect 392 2003 394 2007
rect 398 2003 401 2007
rect 406 2003 408 2007
rect 190 1872 193 1928
rect 290 1888 294 1891
rect 386 1868 390 1871
rect 392 1803 394 1807
rect 398 1803 401 1807
rect 406 1803 408 1807
rect 392 1603 394 1607
rect 398 1603 401 1607
rect 406 1603 408 1607
rect 54 1342 57 1468
rect 78 1442 81 1448
rect 6 1192 9 1298
rect 18 1278 22 1281
rect 14 1242 17 1248
rect 18 1178 22 1181
rect 14 952 17 978
rect 94 612 97 1168
rect 102 782 105 1538
rect 170 1468 174 1471
rect 198 1462 201 1528
rect 422 1522 425 2198
rect 430 1562 433 1918
rect 414 1412 417 1468
rect 392 1403 394 1407
rect 398 1403 401 1407
rect 406 1403 408 1407
rect 110 1272 113 1348
rect 126 1201 129 1348
rect 246 1332 249 1338
rect 122 1198 129 1201
rect 142 1082 145 1278
rect 392 1203 394 1207
rect 398 1203 401 1207
rect 406 1203 408 1207
rect 374 1178 382 1181
rect 374 1142 377 1178
rect 414 1172 417 1198
rect 134 672 137 688
rect 114 628 121 631
rect 118 422 121 628
rect 142 482 145 1078
rect 162 1068 166 1071
rect 150 532 153 928
rect 162 868 166 871
rect 162 738 166 741
rect 182 552 185 1098
rect 118 412 121 418
rect 110 272 113 378
rect 182 362 185 548
rect 210 338 214 341
rect 218 148 222 151
rect 254 142 257 688
rect 270 622 273 1128
rect 294 992 297 1118
rect 392 1003 394 1007
rect 398 1003 401 1007
rect 406 1003 408 1007
rect 374 872 377 928
rect 158 72 161 88
rect 254 72 257 138
rect 286 112 289 618
rect 358 162 361 318
rect 374 182 377 868
rect 392 803 394 807
rect 398 803 401 807
rect 406 803 408 807
rect 386 668 390 671
rect 392 603 394 607
rect 398 603 401 607
rect 406 603 408 607
rect 414 572 417 1058
rect 422 882 425 1118
rect 430 782 433 1558
rect 486 1392 489 2528
rect 494 2122 497 2538
rect 502 2452 505 2578
rect 518 2541 521 2648
rect 514 2538 521 2541
rect 518 2222 521 2538
rect 522 2048 526 2051
rect 526 1912 529 1928
rect 526 1722 529 1908
rect 534 1902 537 2058
rect 534 1872 537 1878
rect 550 1852 553 1878
rect 550 1682 553 1848
rect 510 1462 513 1468
rect 554 1438 561 1441
rect 498 1258 502 1261
rect 446 1248 454 1251
rect 438 582 441 1078
rect 446 562 449 1248
rect 510 1162 513 1318
rect 518 972 521 1438
rect 558 1362 561 1438
rect 526 1262 529 1338
rect 558 1282 561 1358
rect 534 1262 537 1268
rect 566 1202 569 2728
rect 574 2642 577 2738
rect 574 2512 577 2558
rect 574 1732 577 2328
rect 582 2112 585 2488
rect 590 2432 593 2578
rect 606 2552 609 2598
rect 598 2548 606 2551
rect 590 2062 593 2228
rect 590 1802 593 2058
rect 598 1912 601 2548
rect 662 2532 665 2558
rect 614 2448 622 2451
rect 606 1672 609 1718
rect 574 1252 577 1528
rect 530 1008 537 1011
rect 518 852 521 968
rect 534 792 537 1008
rect 542 952 545 1078
rect 392 403 394 407
rect 398 403 401 407
rect 406 403 408 407
rect 382 292 385 348
rect 414 261 417 438
rect 518 282 521 678
rect 534 482 537 788
rect 566 738 574 741
rect 566 532 569 738
rect 582 682 585 1668
rect 614 1542 617 2448
rect 638 2012 641 2158
rect 654 2122 657 2258
rect 646 2092 649 2118
rect 646 2082 649 2088
rect 590 942 593 1518
rect 598 1462 601 1478
rect 606 1452 609 1458
rect 614 1152 617 1498
rect 622 1252 625 1458
rect 630 1271 633 1658
rect 638 1532 641 2008
rect 646 1652 649 2058
rect 650 1468 654 1471
rect 662 1322 665 2528
rect 702 2182 705 2928
rect 726 2822 729 3038
rect 896 2903 898 2907
rect 902 2903 905 2907
rect 910 2903 912 2907
rect 934 2892 937 2968
rect 858 2768 865 2771
rect 726 2322 729 2758
rect 750 2748 758 2751
rect 802 2748 806 2751
rect 750 2572 753 2748
rect 862 2722 865 2768
rect 878 2692 881 2868
rect 1010 2748 1014 2751
rect 886 2692 889 2748
rect 1022 2732 1025 2848
rect 896 2703 898 2707
rect 902 2703 905 2707
rect 910 2703 912 2707
rect 758 2482 761 2548
rect 742 2458 750 2461
rect 742 2312 745 2458
rect 790 2072 793 2298
rect 810 2258 814 2261
rect 798 2072 801 2258
rect 806 2142 809 2158
rect 814 2142 817 2148
rect 670 1972 673 1998
rect 678 1902 681 2048
rect 686 1971 689 2018
rect 702 2002 705 2048
rect 686 1968 694 1971
rect 710 1968 718 1971
rect 710 1932 713 1968
rect 726 1962 729 1968
rect 718 1942 721 1948
rect 686 1542 689 1808
rect 694 1312 697 1418
rect 702 1351 705 1788
rect 710 1642 713 1928
rect 718 1732 721 1778
rect 718 1682 721 1688
rect 710 1432 713 1438
rect 702 1348 710 1351
rect 718 1342 721 1538
rect 726 1462 729 1858
rect 734 1672 737 1768
rect 750 1742 753 2058
rect 770 2048 774 2051
rect 774 2002 777 2028
rect 774 1872 777 1988
rect 782 1962 785 2058
rect 782 1862 785 1958
rect 790 1948 798 1951
rect 766 1572 769 1678
rect 754 1468 758 1471
rect 774 1462 777 1598
rect 630 1268 638 1271
rect 650 1268 657 1271
rect 670 1271 673 1288
rect 666 1268 673 1271
rect 654 1161 657 1268
rect 678 1252 681 1278
rect 686 1162 689 1228
rect 654 1158 665 1161
rect 646 1128 654 1131
rect 646 692 649 1128
rect 662 1062 665 1158
rect 682 1148 689 1151
rect 670 1098 678 1101
rect 662 962 665 1058
rect 670 1042 673 1098
rect 686 1012 689 1148
rect 694 672 697 1188
rect 702 1072 705 1178
rect 718 1142 721 1338
rect 754 1328 758 1331
rect 726 1262 729 1278
rect 702 712 705 838
rect 726 752 729 1258
rect 758 1182 761 1198
rect 766 1162 769 1358
rect 734 792 737 1098
rect 750 1062 753 1148
rect 782 1132 785 1858
rect 790 1842 793 1948
rect 790 1692 793 1838
rect 798 1812 801 1818
rect 806 1732 809 1948
rect 814 1662 817 2018
rect 822 1992 825 2458
rect 830 2262 833 2528
rect 896 2503 898 2507
rect 902 2503 905 2507
rect 910 2503 912 2507
rect 896 2303 898 2307
rect 902 2303 905 2307
rect 910 2303 912 2307
rect 958 2281 961 2328
rect 954 2278 961 2281
rect 842 2258 846 2261
rect 822 1892 825 1918
rect 790 1442 793 1648
rect 814 1571 817 1628
rect 810 1568 817 1571
rect 798 1372 801 1568
rect 814 1502 817 1548
rect 798 1242 801 1368
rect 822 1262 825 1768
rect 830 1482 833 2258
rect 838 2168 846 2171
rect 838 2162 841 2168
rect 842 2148 846 2151
rect 838 1872 841 1888
rect 846 1882 849 1968
rect 854 1801 857 2238
rect 846 1798 857 1801
rect 838 1572 841 1628
rect 846 1591 849 1798
rect 854 1782 857 1788
rect 846 1588 854 1591
rect 862 1552 865 2148
rect 870 2141 873 2168
rect 870 2138 878 2141
rect 870 1902 873 1908
rect 870 1872 873 1878
rect 878 1652 881 2048
rect 886 1752 889 2278
rect 918 2142 921 2148
rect 942 2142 945 2208
rect 966 2182 969 2508
rect 1014 2222 1017 2328
rect 1022 2282 1025 2728
rect 1134 2712 1137 3098
rect 1034 2258 1038 2261
rect 906 2138 910 2141
rect 896 2103 898 2107
rect 902 2103 905 2107
rect 910 2103 912 2107
rect 942 2078 950 2081
rect 934 2032 937 2078
rect 942 2012 945 2078
rect 922 1938 926 1941
rect 896 1903 898 1907
rect 902 1903 905 1907
rect 910 1903 912 1907
rect 914 1828 918 1831
rect 906 1728 910 1731
rect 896 1703 898 1707
rect 902 1703 905 1707
rect 910 1703 912 1707
rect 918 1661 921 1828
rect 966 1732 969 2178
rect 974 1762 977 2218
rect 1010 2168 1017 2171
rect 1014 2142 1017 2168
rect 1046 2102 1049 2698
rect 982 1981 985 2038
rect 982 1978 990 1981
rect 982 1772 985 1978
rect 998 1972 1001 1978
rect 998 1941 1001 1968
rect 994 1938 1001 1941
rect 1006 1872 1009 2088
rect 1002 1858 1006 1861
rect 1014 1732 1017 2028
rect 1022 1962 1025 1978
rect 1022 1938 1030 1941
rect 1022 1722 1025 1938
rect 914 1658 921 1661
rect 838 1522 841 1538
rect 838 1482 841 1498
rect 870 1402 873 1628
rect 878 1532 881 1648
rect 898 1548 902 1551
rect 926 1542 929 1718
rect 838 1241 841 1378
rect 838 1238 846 1241
rect 806 1152 809 1208
rect 742 1058 750 1061
rect 742 812 745 1058
rect 766 1052 769 1078
rect 770 1048 774 1051
rect 766 872 769 898
rect 774 892 777 928
rect 798 881 801 1118
rect 794 878 801 881
rect 754 858 758 861
rect 806 782 809 1148
rect 862 1052 865 1098
rect 870 1092 873 1208
rect 878 1012 881 1528
rect 896 1503 898 1507
rect 902 1503 905 1507
rect 910 1503 912 1507
rect 886 1492 889 1498
rect 886 1342 889 1418
rect 914 1358 918 1361
rect 926 1342 929 1358
rect 922 1318 926 1321
rect 896 1303 898 1307
rect 902 1303 905 1307
rect 910 1303 912 1307
rect 926 1252 929 1268
rect 926 1222 929 1238
rect 926 1192 929 1198
rect 926 1152 929 1158
rect 934 1152 937 1658
rect 950 1582 953 1718
rect 958 1462 961 1658
rect 942 1162 945 1338
rect 958 1302 961 1458
rect 966 1352 969 1718
rect 978 1688 982 1691
rect 974 1312 977 1648
rect 982 1502 985 1568
rect 814 872 817 878
rect 822 852 825 858
rect 734 742 737 778
rect 718 728 726 731
rect 710 462 713 698
rect 718 522 721 728
rect 846 662 849 918
rect 854 902 857 938
rect 886 912 889 1128
rect 896 1103 898 1107
rect 902 1103 905 1107
rect 910 1103 912 1107
rect 934 1082 937 1118
rect 950 1082 953 1248
rect 896 903 898 907
rect 902 903 905 907
rect 910 903 912 907
rect 918 742 921 898
rect 934 801 937 1078
rect 930 798 937 801
rect 534 272 537 278
rect 414 258 422 261
rect 392 203 394 207
rect 398 203 401 207
rect 406 203 408 207
rect 478 82 481 268
rect 494 142 497 168
rect 358 11 361 78
rect 542 22 545 288
rect 550 92 553 388
rect 550 62 553 68
rect 558 22 561 438
rect 354 8 361 11
rect 574 11 577 98
rect 570 8 577 11
rect 630 11 633 268
rect 678 222 681 418
rect 710 352 713 458
rect 770 398 774 401
rect 790 392 793 438
rect 854 422 857 728
rect 896 703 898 707
rect 902 703 905 707
rect 910 703 912 707
rect 918 692 921 698
rect 942 672 945 908
rect 958 552 961 1298
rect 974 1132 977 1268
rect 982 1202 985 1498
rect 1014 1342 1017 1668
rect 1030 1472 1033 1878
rect 1046 1372 1049 1738
rect 1054 1322 1057 2168
rect 1062 2112 1065 2338
rect 1070 2062 1073 2448
rect 1078 2082 1081 2308
rect 1074 2058 1078 2061
rect 1070 1762 1073 1858
rect 1074 1728 1081 1731
rect 1062 1352 1065 1728
rect 1078 1652 1081 1728
rect 1086 1592 1089 2318
rect 1094 2302 1097 2448
rect 1134 2382 1137 2538
rect 1118 2261 1121 2338
rect 1142 2332 1145 2368
rect 1118 2258 1126 2261
rect 1118 2022 1121 2258
rect 1102 1682 1105 2008
rect 1142 1982 1145 2028
rect 1138 1958 1142 1961
rect 1114 1908 1121 1911
rect 1118 1892 1121 1908
rect 1134 1902 1137 1938
rect 1142 1932 1145 1938
rect 1126 1762 1129 1878
rect 1134 1872 1137 1878
rect 1134 1692 1137 1798
rect 1142 1722 1145 1908
rect 1150 1761 1153 2158
rect 1158 2051 1161 2318
rect 1166 2132 1169 2738
rect 1174 2122 1177 3098
rect 1202 2868 1209 2871
rect 1206 2702 1209 2868
rect 1182 2212 1185 2648
rect 1158 2048 1166 2051
rect 1174 2042 1177 2048
rect 1158 1942 1161 1998
rect 1150 1758 1158 1761
rect 1166 1722 1169 1958
rect 1138 1668 1142 1671
rect 1122 1648 1126 1651
rect 982 1142 985 1198
rect 966 1062 969 1108
rect 982 1062 985 1068
rect 990 882 993 1068
rect 974 842 977 848
rect 722 318 726 321
rect 782 312 785 388
rect 886 342 889 518
rect 896 503 898 507
rect 902 503 905 507
rect 910 503 912 507
rect 918 412 921 508
rect 974 352 977 548
rect 982 382 985 748
rect 998 512 1001 1068
rect 1006 942 1009 1318
rect 1014 872 1017 1298
rect 1070 1272 1073 1288
rect 1046 1092 1049 1118
rect 1030 1018 1038 1021
rect 1022 642 1025 898
rect 1030 672 1033 1018
rect 1038 982 1041 1008
rect 1046 942 1049 1068
rect 1054 952 1057 1238
rect 1078 1212 1081 1518
rect 1094 1292 1097 1508
rect 1102 1482 1105 1648
rect 1106 1288 1110 1291
rect 1062 1022 1065 1158
rect 1070 1152 1073 1158
rect 1038 862 1041 918
rect 1070 742 1073 1068
rect 1078 1062 1081 1068
rect 1086 942 1089 1278
rect 1094 932 1097 1168
rect 1102 1162 1105 1178
rect 1110 961 1113 1218
rect 1118 1192 1121 1588
rect 1126 1281 1129 1548
rect 1134 1342 1137 1528
rect 1126 1278 1134 1281
rect 1126 1162 1129 1278
rect 1106 958 1113 961
rect 1078 642 1081 698
rect 1078 592 1081 638
rect 1094 562 1097 688
rect 1102 542 1105 698
rect 1110 542 1113 888
rect 1118 822 1121 1148
rect 1134 1002 1137 1258
rect 1142 1222 1145 1458
rect 1166 1342 1169 1668
rect 1174 1352 1177 1968
rect 1182 1262 1185 2178
rect 1190 1642 1193 2598
rect 1214 2402 1217 2648
rect 1238 2492 1241 2668
rect 1246 2622 1249 2918
rect 1254 2712 1257 2868
rect 1270 2742 1273 2818
rect 1262 2738 1270 2741
rect 1198 2052 1201 2268
rect 1206 1862 1209 2268
rect 1230 2132 1233 2488
rect 1242 1938 1246 1941
rect 1254 1931 1257 2318
rect 1246 1928 1257 1931
rect 1206 1682 1209 1788
rect 1230 1742 1233 1808
rect 1246 1732 1249 1928
rect 1262 1801 1265 2738
rect 1286 2222 1289 2628
rect 1302 2272 1305 2638
rect 1310 2232 1313 2248
rect 1286 2062 1289 2218
rect 1278 1942 1281 1968
rect 1254 1798 1265 1801
rect 1270 1802 1273 1938
rect 1286 1862 1289 1878
rect 1294 1862 1297 2108
rect 1302 1932 1305 2138
rect 1326 2082 1329 2808
rect 1334 2282 1337 3098
rect 1416 3003 1418 3007
rect 1422 3003 1425 3007
rect 1430 3003 1432 3007
rect 1462 2952 1465 2958
rect 1470 2852 1473 3088
rect 1602 3058 1609 3061
rect 1478 2968 1486 2971
rect 1478 2892 1481 2968
rect 1566 2922 1569 3028
rect 1558 2862 1561 2868
rect 1416 2803 1418 2807
rect 1422 2803 1425 2807
rect 1430 2803 1432 2807
rect 1370 2458 1374 2461
rect 1354 2448 1358 2451
rect 1318 1992 1321 2028
rect 1198 1678 1206 1681
rect 1150 1238 1158 1241
rect 1142 1032 1145 1148
rect 1150 1052 1153 1238
rect 1166 1012 1169 1258
rect 1166 972 1169 1008
rect 1154 948 1158 951
rect 1134 942 1137 948
rect 1126 761 1129 908
rect 1142 882 1145 948
rect 1122 758 1129 761
rect 1126 602 1129 748
rect 1134 742 1137 758
rect 1062 338 1070 341
rect 896 303 898 307
rect 902 303 905 307
rect 910 303 912 307
rect 918 272 921 308
rect 950 292 953 298
rect 838 232 841 248
rect 694 142 697 158
rect 974 152 977 168
rect 990 152 993 158
rect 896 103 898 107
rect 902 103 905 107
rect 910 103 912 107
rect 630 8 638 11
rect 774 11 777 98
rect 770 8 777 11
rect 1006 11 1009 298
rect 1062 272 1065 338
rect 1110 282 1113 538
rect 1118 432 1121 598
rect 1134 452 1137 508
rect 1142 471 1145 868
rect 1142 468 1150 471
rect 1174 422 1177 1058
rect 1182 962 1185 1178
rect 1190 752 1193 1488
rect 1198 1152 1201 1678
rect 1214 1362 1217 1648
rect 1238 1522 1241 1718
rect 1254 1462 1257 1798
rect 1286 1772 1289 1858
rect 1278 1681 1281 1688
rect 1302 1682 1305 1728
rect 1278 1678 1286 1681
rect 1262 1542 1265 1628
rect 1262 1528 1265 1538
rect 1206 1282 1209 1298
rect 1206 1132 1209 1138
rect 1206 1112 1209 1118
rect 1198 432 1201 978
rect 1206 952 1209 958
rect 1214 922 1217 1358
rect 1222 962 1225 1368
rect 1230 1332 1233 1338
rect 1230 1142 1233 1168
rect 1234 1128 1238 1131
rect 1222 952 1225 958
rect 1230 942 1233 948
rect 1234 668 1241 671
rect 1226 648 1233 651
rect 1150 322 1153 328
rect 1118 162 1121 218
rect 1182 162 1185 358
rect 1206 332 1209 628
rect 1214 332 1217 528
rect 1222 482 1225 488
rect 1230 412 1233 648
rect 1238 532 1241 668
rect 1246 522 1249 1118
rect 1254 972 1257 1458
rect 1274 1348 1278 1351
rect 1302 1342 1305 1408
rect 1262 1112 1265 1338
rect 1310 1322 1313 1968
rect 1326 1932 1329 2078
rect 1318 1822 1321 1878
rect 1318 1682 1321 1808
rect 1326 1752 1329 1908
rect 1334 1702 1337 2268
rect 1342 1832 1345 2358
rect 1382 2352 1385 2588
rect 1350 1942 1353 2098
rect 1326 1362 1329 1368
rect 1334 1362 1337 1618
rect 1342 1382 1345 1818
rect 1350 1361 1353 1798
rect 1358 1562 1361 2208
rect 1382 2152 1385 2348
rect 1390 2342 1393 2478
rect 1398 2402 1401 2678
rect 1416 2603 1418 2607
rect 1422 2603 1425 2607
rect 1430 2603 1432 2607
rect 1438 2502 1441 2808
rect 1510 2532 1513 2538
rect 1446 2452 1449 2498
rect 1514 2408 1518 2411
rect 1416 2403 1418 2407
rect 1422 2403 1425 2407
rect 1430 2403 1432 2407
rect 1398 2342 1401 2348
rect 1366 1952 1369 1968
rect 1366 1732 1369 1938
rect 1382 1912 1385 1948
rect 1374 1842 1377 1848
rect 1378 1748 1382 1751
rect 1386 1718 1390 1721
rect 1366 1662 1369 1668
rect 1382 1662 1385 1688
rect 1366 1572 1369 1648
rect 1374 1542 1377 1658
rect 1350 1358 1358 1361
rect 1350 1342 1353 1358
rect 1342 1271 1345 1308
rect 1338 1268 1345 1271
rect 1290 1258 1294 1261
rect 1326 1252 1329 1268
rect 1334 1152 1337 1258
rect 1270 1082 1273 1098
rect 1266 1078 1270 1081
rect 1278 1072 1281 1128
rect 1254 952 1257 968
rect 1266 948 1270 951
rect 1278 862 1281 1068
rect 1302 1062 1305 1068
rect 1286 912 1289 958
rect 1310 802 1313 1058
rect 1318 862 1321 978
rect 1326 962 1329 1148
rect 1334 932 1337 1088
rect 1342 972 1345 1258
rect 1350 1122 1353 1288
rect 1358 1172 1361 1218
rect 1342 922 1345 968
rect 1350 962 1353 1078
rect 1358 922 1361 1158
rect 1366 952 1369 1468
rect 1374 1352 1377 1358
rect 1374 1282 1377 1338
rect 1390 1322 1393 1488
rect 1382 1292 1385 1298
rect 1382 1202 1385 1278
rect 1390 1192 1393 1308
rect 1374 1112 1377 1148
rect 1362 918 1369 921
rect 1326 702 1329 918
rect 1334 742 1337 898
rect 1254 652 1257 668
rect 1310 651 1313 678
rect 1310 648 1318 651
rect 1230 402 1233 408
rect 1230 272 1233 388
rect 1238 342 1241 488
rect 1254 481 1257 518
rect 1270 482 1273 558
rect 1278 548 1286 551
rect 1254 478 1262 481
rect 1278 352 1281 548
rect 1238 318 1246 321
rect 1198 192 1201 268
rect 1114 138 1118 141
rect 1150 141 1153 148
rect 1150 138 1158 141
rect 1022 52 1025 88
rect 1030 72 1033 138
rect 1090 128 1094 131
rect 1038 82 1041 128
rect 1102 72 1105 78
rect 1006 8 1014 11
rect 1198 11 1201 188
rect 1214 172 1217 198
rect 1230 52 1233 248
rect 1238 72 1241 318
rect 1266 298 1270 301
rect 1246 162 1249 258
rect 1254 142 1257 148
rect 1262 132 1265 178
rect 1274 158 1278 161
rect 1286 112 1289 538
rect 1298 478 1302 481
rect 1310 352 1313 368
rect 1294 332 1297 338
rect 1350 322 1353 838
rect 1366 832 1369 918
rect 1366 742 1369 748
rect 1366 462 1369 608
rect 1358 418 1366 421
rect 1306 188 1310 191
rect 1314 138 1318 141
rect 1250 78 1254 81
rect 1326 72 1329 238
rect 1334 122 1337 318
rect 1350 262 1353 318
rect 1342 92 1345 118
rect 1358 92 1361 418
rect 1374 161 1377 1008
rect 1382 852 1385 1138
rect 1398 1132 1401 2268
rect 1406 2072 1409 2388
rect 1416 2203 1418 2207
rect 1422 2203 1425 2207
rect 1430 2203 1432 2207
rect 1438 2162 1441 2298
rect 1518 2102 1521 2338
rect 1526 2132 1529 2158
rect 1534 2112 1537 2668
rect 1542 2582 1545 2678
rect 1406 1642 1409 2068
rect 1416 2003 1418 2007
rect 1422 2003 1425 2007
rect 1430 2003 1432 2007
rect 1458 1978 1462 1981
rect 1414 1842 1417 1928
rect 1416 1803 1418 1807
rect 1422 1803 1425 1807
rect 1430 1803 1432 1807
rect 1438 1672 1441 1928
rect 1446 1922 1449 1938
rect 1462 1892 1465 1898
rect 1470 1892 1473 2068
rect 1482 1928 1489 1931
rect 1454 1832 1457 1838
rect 1446 1672 1449 1678
rect 1454 1662 1457 1828
rect 1462 1642 1465 1858
rect 1406 1592 1409 1608
rect 1416 1603 1418 1607
rect 1422 1603 1425 1607
rect 1430 1603 1432 1607
rect 1462 1602 1465 1638
rect 1462 1552 1465 1558
rect 1406 1462 1409 1508
rect 1390 902 1393 1108
rect 1398 902 1401 1118
rect 1406 1072 1409 1438
rect 1438 1412 1441 1538
rect 1416 1403 1418 1407
rect 1422 1403 1425 1407
rect 1430 1403 1432 1407
rect 1446 1352 1449 1538
rect 1414 1332 1417 1348
rect 1418 1258 1422 1261
rect 1416 1203 1418 1207
rect 1422 1203 1425 1207
rect 1430 1203 1432 1207
rect 1438 1191 1441 1208
rect 1430 1188 1441 1191
rect 1430 1182 1433 1188
rect 1416 1003 1418 1007
rect 1422 1003 1425 1007
rect 1430 1003 1432 1007
rect 1394 888 1398 891
rect 1398 822 1401 868
rect 1382 412 1385 818
rect 1398 662 1401 818
rect 1406 652 1409 808
rect 1416 803 1418 807
rect 1422 803 1425 807
rect 1430 803 1432 807
rect 1422 712 1425 768
rect 1430 752 1433 778
rect 1438 732 1441 958
rect 1416 603 1418 607
rect 1422 603 1425 607
rect 1430 603 1432 607
rect 1438 582 1441 718
rect 1446 682 1449 938
rect 1454 872 1457 1448
rect 1462 1382 1465 1498
rect 1470 1452 1473 1848
rect 1478 1552 1481 1838
rect 1486 1762 1489 1928
rect 1462 1062 1465 1358
rect 1470 1272 1473 1398
rect 1478 1342 1481 1538
rect 1486 1372 1489 1748
rect 1494 1652 1497 2038
rect 1494 1482 1497 1578
rect 1502 1562 1505 1918
rect 1510 1872 1513 1878
rect 1510 1752 1513 1758
rect 1510 1652 1513 1658
rect 1494 1472 1497 1478
rect 1502 1442 1505 1458
rect 1494 1382 1497 1388
rect 1486 1352 1489 1368
rect 1510 1342 1513 1548
rect 1518 1522 1521 2038
rect 1542 1972 1545 2108
rect 1526 1732 1529 1878
rect 1534 1722 1537 1848
rect 1526 1672 1529 1708
rect 1534 1482 1537 1628
rect 1542 1602 1545 1768
rect 1550 1632 1553 2518
rect 1558 1822 1561 1998
rect 1574 1962 1577 2228
rect 1598 2132 1601 2888
rect 1606 2272 1609 3058
rect 1674 2948 1678 2951
rect 1694 2912 1697 3098
rect 1750 2872 1753 2878
rect 1614 2572 1617 2718
rect 1614 2332 1617 2568
rect 1622 2492 1625 2738
rect 1630 2342 1633 2528
rect 1662 2462 1665 2668
rect 1694 2492 1697 2608
rect 1682 2478 1686 2481
rect 1646 2438 1654 2441
rect 1622 2322 1625 2328
rect 1638 2252 1641 2408
rect 1646 2392 1649 2438
rect 1646 2282 1649 2388
rect 1630 2248 1638 2251
rect 1582 1952 1585 2038
rect 1582 1932 1585 1948
rect 1598 1912 1601 2128
rect 1606 1972 1609 2118
rect 1614 1932 1617 1998
rect 1574 1891 1577 1898
rect 1570 1888 1577 1891
rect 1574 1712 1577 1718
rect 1582 1632 1585 1728
rect 1606 1662 1609 1668
rect 1550 1532 1553 1548
rect 1470 1142 1473 1258
rect 1462 1032 1465 1058
rect 1470 1052 1473 1098
rect 1478 1082 1481 1338
rect 1486 1322 1489 1328
rect 1486 1102 1489 1308
rect 1494 1232 1497 1248
rect 1494 1192 1497 1208
rect 1478 1058 1486 1061
rect 1466 1018 1473 1021
rect 1470 892 1473 1018
rect 1454 842 1457 848
rect 1366 158 1377 161
rect 1390 222 1393 518
rect 1330 28 1334 31
rect 1194 8 1201 11
rect 1366 12 1369 158
rect 1374 132 1377 148
rect 1374 72 1377 128
rect 1390 122 1393 218
rect 1382 62 1385 98
rect 1398 92 1401 188
rect 1406 171 1409 568
rect 1418 548 1422 551
rect 1446 542 1449 678
rect 1446 472 1449 478
rect 1454 472 1457 748
rect 1462 742 1465 888
rect 1462 712 1465 738
rect 1462 672 1465 698
rect 1462 562 1465 568
rect 1416 403 1418 407
rect 1422 403 1425 407
rect 1430 403 1432 407
rect 1470 302 1473 718
rect 1478 652 1481 1058
rect 1486 741 1489 988
rect 1494 942 1497 1128
rect 1502 912 1505 1248
rect 1510 1152 1513 1308
rect 1510 992 1513 1138
rect 1518 992 1521 1478
rect 1526 1322 1529 1378
rect 1550 1342 1553 1528
rect 1526 1262 1529 1318
rect 1542 1282 1545 1298
rect 1534 1232 1537 1258
rect 1542 1242 1545 1248
rect 1550 1202 1553 1308
rect 1558 1162 1561 1498
rect 1566 1422 1569 1458
rect 1574 1332 1577 1348
rect 1582 1342 1585 1528
rect 1606 1522 1609 1528
rect 1590 1452 1593 1458
rect 1614 1362 1617 1898
rect 1622 1512 1625 2178
rect 1630 1882 1633 2248
rect 1638 2052 1641 2058
rect 1654 1912 1657 2428
rect 1662 2292 1665 2318
rect 1670 2312 1673 2468
rect 1682 2458 1686 2461
rect 1702 2392 1705 2438
rect 1670 2282 1673 2308
rect 1670 1872 1673 2278
rect 1678 2212 1681 2288
rect 1686 2252 1689 2348
rect 1698 2278 1702 2281
rect 1662 1852 1665 1868
rect 1638 1602 1641 1838
rect 1686 1802 1689 2248
rect 1694 2092 1697 2098
rect 1694 1862 1697 2068
rect 1666 1758 1670 1761
rect 1654 1682 1657 1698
rect 1646 1592 1649 1608
rect 1634 1568 1638 1571
rect 1654 1562 1657 1598
rect 1662 1592 1665 1748
rect 1678 1652 1681 1718
rect 1686 1672 1689 1798
rect 1702 1732 1705 2118
rect 1710 2082 1713 2758
rect 1750 2552 1753 2588
rect 1734 2482 1737 2488
rect 1718 2262 1721 2278
rect 1734 2162 1737 2258
rect 1718 1882 1721 2078
rect 1726 2062 1729 2068
rect 1734 1942 1737 2158
rect 1750 1992 1753 2448
rect 1758 2312 1761 2358
rect 1766 2352 1769 2678
rect 1798 2442 1801 2738
rect 1814 2552 1817 2558
rect 1806 2532 1809 2538
rect 1786 2348 1790 2351
rect 1774 2232 1777 2278
rect 1806 2252 1809 2488
rect 1750 1972 1753 1988
rect 1750 1952 1753 1958
rect 1758 1922 1761 2178
rect 1766 2162 1769 2168
rect 1766 1882 1769 1888
rect 1722 1868 1726 1871
rect 1746 1858 1750 1861
rect 1654 1552 1657 1558
rect 1662 1552 1665 1588
rect 1678 1542 1681 1648
rect 1574 1322 1577 1328
rect 1566 1232 1569 1308
rect 1534 1122 1537 1128
rect 1530 1088 1534 1091
rect 1542 1072 1545 1078
rect 1510 962 1513 968
rect 1518 912 1521 988
rect 1550 922 1553 1128
rect 1558 962 1561 1128
rect 1566 1082 1569 1088
rect 1566 1042 1569 1058
rect 1574 1022 1577 1178
rect 1582 1082 1585 1338
rect 1590 1282 1593 1308
rect 1598 1272 1601 1348
rect 1610 1318 1614 1321
rect 1622 1282 1625 1498
rect 1678 1492 1681 1518
rect 1686 1482 1689 1508
rect 1638 1382 1641 1448
rect 1646 1412 1649 1448
rect 1634 1358 1638 1361
rect 1634 1318 1641 1321
rect 1638 1312 1641 1318
rect 1606 1222 1609 1278
rect 1630 1252 1633 1268
rect 1582 1022 1585 1048
rect 1558 912 1561 918
rect 1534 908 1542 911
rect 1494 802 1497 808
rect 1486 738 1494 741
rect 1486 662 1489 668
rect 1442 268 1446 271
rect 1478 242 1481 538
rect 1486 392 1489 478
rect 1494 472 1497 738
rect 1510 662 1513 878
rect 1518 542 1521 668
rect 1534 462 1537 908
rect 1486 262 1489 268
rect 1494 262 1497 368
rect 1518 362 1521 458
rect 1478 232 1481 238
rect 1416 203 1418 207
rect 1422 203 1425 207
rect 1430 203 1432 207
rect 1406 168 1417 171
rect 1406 142 1409 148
rect 1414 132 1417 168
rect 1438 82 1441 208
rect 1510 82 1513 228
rect 1518 102 1521 268
rect 1526 222 1529 458
rect 1550 442 1553 788
rect 1558 622 1561 698
rect 1566 652 1569 938
rect 1574 632 1577 918
rect 1582 842 1585 998
rect 1590 842 1593 1048
rect 1558 532 1561 618
rect 1582 492 1585 708
rect 1566 468 1574 471
rect 1542 362 1545 428
rect 1550 152 1553 338
rect 1566 162 1569 468
rect 1590 362 1593 798
rect 1598 782 1601 1198
rect 1606 932 1609 1218
rect 1622 1122 1625 1128
rect 1622 1112 1625 1118
rect 1630 1092 1633 1178
rect 1598 602 1601 678
rect 1606 662 1609 928
rect 1622 882 1625 1068
rect 1638 1062 1641 1248
rect 1646 1062 1649 1378
rect 1654 1242 1657 1408
rect 1662 1222 1665 1448
rect 1674 1438 1678 1441
rect 1674 1348 1678 1351
rect 1654 1042 1657 1118
rect 1662 1092 1665 1158
rect 1670 1118 1678 1121
rect 1638 922 1641 1028
rect 1654 992 1657 1038
rect 1650 928 1654 931
rect 1654 842 1657 868
rect 1670 842 1673 1118
rect 1686 1062 1689 1458
rect 1694 1322 1697 1658
rect 1682 1048 1689 1051
rect 1686 982 1689 1048
rect 1686 882 1689 898
rect 1686 871 1689 878
rect 1682 868 1689 871
rect 1670 832 1673 838
rect 1614 722 1617 728
rect 1614 682 1617 708
rect 1614 658 1622 661
rect 1614 522 1617 658
rect 1638 572 1641 808
rect 1646 722 1649 798
rect 1694 752 1697 1148
rect 1702 1122 1705 1668
rect 1718 1572 1721 1738
rect 1758 1642 1761 1858
rect 1774 1782 1777 1988
rect 1782 1652 1785 2238
rect 1794 2228 1798 2231
rect 1806 1942 1809 2148
rect 1806 1912 1809 1938
rect 1802 1718 1806 1721
rect 1790 1712 1793 1718
rect 1794 1708 1801 1711
rect 1798 1692 1801 1708
rect 1710 1242 1713 1478
rect 1718 1392 1721 1568
rect 1738 1558 1742 1561
rect 1726 1472 1729 1508
rect 1758 1482 1761 1528
rect 1758 1472 1761 1478
rect 1774 1472 1777 1648
rect 1790 1512 1793 1688
rect 1798 1542 1801 1688
rect 1806 1672 1809 1688
rect 1782 1452 1785 1488
rect 1794 1448 1798 1451
rect 1726 1382 1729 1398
rect 1734 1332 1737 1348
rect 1718 1312 1721 1328
rect 1730 1318 1734 1321
rect 1750 1321 1753 1388
rect 1758 1362 1761 1428
rect 1746 1318 1753 1321
rect 1742 1232 1745 1278
rect 1758 1272 1761 1348
rect 1766 1322 1769 1328
rect 1758 1252 1761 1258
rect 1750 1242 1753 1248
rect 1766 1232 1769 1258
rect 1750 1222 1753 1228
rect 1718 1152 1721 1168
rect 1702 1072 1705 1118
rect 1710 1062 1713 1118
rect 1726 1062 1729 1158
rect 1710 1012 1713 1058
rect 1746 958 1750 961
rect 1758 952 1761 1168
rect 1774 1102 1777 1348
rect 1798 1262 1801 1318
rect 1766 1072 1769 1078
rect 1774 1072 1777 1088
rect 1702 841 1705 928
rect 1722 888 1726 891
rect 1722 878 1726 881
rect 1730 868 1734 871
rect 1702 838 1710 841
rect 1702 802 1705 808
rect 1702 742 1705 748
rect 1662 721 1665 728
rect 1658 718 1665 721
rect 1654 708 1662 711
rect 1606 282 1609 478
rect 1646 402 1649 708
rect 1550 142 1553 148
rect 1502 72 1505 78
rect 1566 62 1569 158
rect 1590 92 1593 278
rect 1598 52 1601 248
rect 1606 202 1609 278
rect 1610 148 1614 151
rect 1642 138 1646 141
rect 1654 122 1657 708
rect 1694 702 1697 718
rect 1674 658 1681 661
rect 1662 552 1665 578
rect 1678 532 1681 658
rect 1702 492 1705 738
rect 1710 642 1713 838
rect 1718 762 1721 868
rect 1718 742 1721 758
rect 1734 592 1737 748
rect 1742 502 1745 748
rect 1758 652 1761 928
rect 1766 868 1774 871
rect 1766 652 1769 868
rect 1782 832 1785 1218
rect 1790 992 1793 1178
rect 1806 1052 1809 1628
rect 1814 1622 1817 2378
rect 1822 2332 1825 2788
rect 1830 2422 1833 2908
rect 1830 2342 1833 2368
rect 1838 2092 1841 2458
rect 1846 2432 1849 3058
rect 1858 2528 1862 2531
rect 1870 2521 1873 2668
rect 1862 2518 1873 2521
rect 1854 2462 1857 2468
rect 1846 2342 1849 2398
rect 1862 2342 1865 2518
rect 1862 2312 1865 2318
rect 1846 2262 1849 2308
rect 1814 1552 1817 1558
rect 1822 1402 1825 2048
rect 1834 2008 1838 2011
rect 1854 1992 1857 2288
rect 1862 2252 1865 2298
rect 1870 2262 1873 2468
rect 1866 2038 1870 2041
rect 1850 1908 1857 1911
rect 1838 1772 1841 1838
rect 1854 1822 1857 1908
rect 1838 1622 1841 1768
rect 1822 1282 1825 1308
rect 1822 1192 1825 1228
rect 1822 1131 1825 1188
rect 1818 1128 1825 1131
rect 1822 1092 1825 1108
rect 1790 952 1793 988
rect 1802 878 1809 881
rect 1794 838 1801 841
rect 1798 792 1801 838
rect 1806 812 1809 878
rect 1802 738 1809 741
rect 1806 722 1809 738
rect 1814 722 1817 1068
rect 1822 942 1825 1088
rect 1830 1052 1833 1538
rect 1838 1432 1841 1538
rect 1826 878 1830 881
rect 1838 732 1841 1358
rect 1846 882 1849 1728
rect 1854 1182 1857 1768
rect 1862 1222 1865 1638
rect 1870 1622 1873 1988
rect 1878 1882 1881 2918
rect 1886 2102 1889 2858
rect 1902 2812 1905 3098
rect 1910 2772 1913 3098
rect 1928 2903 1930 2907
rect 1934 2903 1937 2907
rect 1942 2903 1944 2907
rect 1918 2712 1921 2778
rect 1928 2703 1930 2707
rect 1934 2703 1937 2707
rect 1942 2703 1944 2707
rect 1894 2342 1897 2638
rect 1918 2482 1921 2538
rect 1928 2503 1930 2507
rect 1934 2503 1937 2507
rect 1942 2503 1944 2507
rect 1950 2492 1953 2498
rect 1886 2012 1889 2018
rect 1878 1782 1881 1878
rect 1894 1862 1897 2338
rect 1902 2242 1905 2438
rect 1902 2032 1905 2148
rect 1910 2112 1913 2448
rect 1918 1942 1921 2478
rect 1928 2303 1930 2307
rect 1934 2303 1937 2307
rect 1942 2303 1944 2307
rect 1928 2103 1930 2107
rect 1934 2103 1937 2107
rect 1942 2103 1944 2107
rect 1934 1972 1937 2048
rect 1950 2042 1953 2388
rect 1958 2372 1961 3018
rect 1982 2822 1985 2908
rect 1966 2292 1969 2548
rect 1974 2102 1977 2368
rect 1982 2362 1985 2658
rect 1998 2542 2001 2808
rect 2046 2682 2049 2968
rect 2054 2682 2057 2738
rect 2046 2602 2049 2618
rect 2014 2562 2017 2568
rect 1998 2412 2001 2538
rect 1982 2302 1985 2358
rect 1994 2338 1998 2341
rect 2006 2262 2009 2498
rect 2014 2302 2017 2558
rect 2054 2462 2057 2628
rect 2062 2542 2065 2798
rect 2054 2442 2057 2458
rect 2062 2362 2065 2378
rect 2014 2262 2017 2278
rect 1986 2248 1990 2251
rect 2026 2248 2030 2251
rect 2006 2242 2009 2248
rect 1986 2228 1990 2231
rect 2006 2182 2009 2198
rect 2006 2142 2009 2178
rect 1998 2132 2001 2138
rect 2014 2132 2017 2238
rect 1966 2022 1969 2048
rect 1946 1988 1950 1991
rect 1966 1982 1969 2018
rect 1902 1938 1910 1941
rect 1934 1932 1937 1948
rect 2022 1941 2025 2198
rect 2030 2012 2033 2158
rect 2018 1938 2025 1941
rect 2038 1952 2041 2338
rect 2058 2168 2062 2171
rect 2062 2032 2065 2128
rect 2070 1972 2073 2588
rect 2086 2582 2089 2748
rect 2094 2692 2097 2768
rect 2094 2532 2097 2648
rect 2090 2528 2094 2531
rect 2086 2462 2089 2478
rect 2086 2451 2089 2458
rect 2082 2448 2089 2451
rect 2110 2432 2113 2748
rect 2142 2731 2145 3088
rect 2158 2882 2161 2898
rect 2154 2858 2161 2861
rect 2158 2732 2161 2858
rect 2142 2728 2150 2731
rect 2078 2352 2081 2368
rect 2094 2342 2097 2348
rect 2086 2062 2089 2328
rect 2110 2092 2113 2298
rect 2118 2172 2121 2458
rect 2142 2412 2145 2728
rect 2134 2312 2137 2328
rect 2130 2258 2134 2261
rect 1886 1702 1889 1718
rect 1870 1442 1873 1568
rect 1886 1522 1889 1578
rect 1894 1552 1897 1808
rect 1886 1482 1889 1518
rect 1894 1502 1897 1548
rect 1894 1472 1897 1478
rect 1870 1322 1873 1368
rect 1882 1358 1886 1361
rect 1890 1348 1897 1351
rect 1882 1318 1889 1321
rect 1886 1282 1889 1318
rect 1862 1082 1865 1138
rect 1854 1072 1857 1078
rect 1854 1062 1857 1068
rect 1854 942 1857 968
rect 1854 822 1857 928
rect 1862 832 1865 1068
rect 1870 1042 1873 1128
rect 1870 952 1873 1038
rect 1886 1032 1889 1278
rect 1894 1272 1897 1348
rect 1870 892 1873 918
rect 1862 802 1865 808
rect 1834 718 1841 721
rect 1778 688 1782 691
rect 1806 552 1809 718
rect 1702 402 1705 488
rect 1742 402 1745 498
rect 1758 472 1761 528
rect 1678 302 1681 348
rect 1726 342 1729 348
rect 1670 92 1673 298
rect 1718 142 1721 248
rect 1710 132 1713 138
rect 1726 132 1729 338
rect 1758 312 1761 468
rect 1774 462 1777 508
rect 1782 322 1785 528
rect 1838 452 1841 718
rect 1846 692 1849 698
rect 1870 682 1873 808
rect 1878 682 1881 1008
rect 1886 912 1889 918
rect 1858 568 1862 571
rect 1878 412 1881 648
rect 1798 372 1801 378
rect 1782 282 1785 318
rect 1806 112 1809 378
rect 1886 342 1889 878
rect 1894 672 1897 1188
rect 1902 842 1905 1898
rect 1918 1882 1921 1908
rect 1928 1903 1930 1907
rect 1934 1903 1937 1907
rect 1942 1903 1944 1907
rect 1990 1762 1993 1778
rect 1974 1732 1977 1738
rect 2006 1732 2009 1858
rect 2014 1742 2017 1938
rect 1958 1712 1961 1728
rect 1928 1703 1930 1707
rect 1934 1703 1937 1707
rect 1942 1703 1944 1707
rect 1926 1672 1929 1688
rect 1914 1648 1921 1651
rect 1918 1642 1921 1648
rect 1970 1628 1974 1631
rect 1910 1482 1913 1508
rect 1910 1432 1913 1438
rect 1918 1392 1921 1618
rect 1966 1602 1969 1618
rect 1926 1532 1929 1538
rect 1928 1503 1930 1507
rect 1934 1503 1937 1507
rect 1942 1503 1944 1507
rect 1926 1422 1929 1438
rect 1942 1382 1945 1458
rect 1910 1312 1913 1338
rect 1928 1303 1930 1307
rect 1934 1303 1937 1307
rect 1942 1303 1944 1307
rect 1902 712 1905 828
rect 1910 812 1913 1228
rect 1918 1162 1921 1178
rect 1918 1002 1921 1118
rect 1928 1103 1930 1107
rect 1934 1103 1937 1107
rect 1942 1103 1944 1107
rect 1950 1072 1953 1258
rect 1958 1172 1961 1538
rect 1966 1362 1969 1588
rect 1974 1522 1977 1558
rect 1974 1331 1977 1508
rect 1966 1328 1977 1331
rect 1958 1061 1961 1128
rect 1950 1058 1961 1061
rect 1942 932 1945 1018
rect 1902 632 1905 708
rect 1918 382 1921 928
rect 1928 903 1930 907
rect 1934 903 1937 907
rect 1942 903 1944 907
rect 1938 848 1942 851
rect 1950 732 1953 1058
rect 1928 703 1930 707
rect 1934 703 1937 707
rect 1942 703 1944 707
rect 1926 622 1929 678
rect 1958 662 1961 1008
rect 1966 752 1969 1328
rect 1982 1242 1985 1728
rect 2006 1672 2009 1698
rect 2014 1672 2017 1678
rect 2038 1662 2041 1948
rect 2054 1852 2057 1888
rect 2066 1858 2070 1861
rect 2054 1782 2057 1798
rect 2046 1752 2049 1758
rect 2062 1751 2065 1758
rect 2058 1748 2065 1751
rect 2062 1742 2065 1748
rect 2046 1702 2049 1738
rect 2006 1642 2009 1648
rect 2070 1622 2073 1818
rect 2078 1772 2081 1908
rect 2086 1772 2089 1878
rect 2102 1852 2105 1858
rect 2082 1608 2086 1611
rect 1990 1532 1993 1598
rect 2002 1558 2006 1561
rect 2094 1542 2097 1848
rect 2102 1742 2105 1808
rect 2102 1722 2105 1738
rect 2102 1542 2105 1658
rect 2110 1642 2113 2088
rect 2142 1962 2145 1978
rect 2118 1612 2121 1958
rect 2010 1448 2014 1451
rect 1974 1182 1977 1198
rect 1974 1082 1977 1178
rect 1990 992 1993 1438
rect 2002 1388 2006 1391
rect 2114 1378 2118 1381
rect 2006 1358 2014 1361
rect 2006 1352 2009 1358
rect 2014 1282 2017 1308
rect 2038 1282 2041 1288
rect 1998 1152 2001 1218
rect 2002 1128 2006 1131
rect 1990 922 1993 968
rect 1974 918 1982 921
rect 1974 872 1977 918
rect 1974 592 1977 838
rect 1990 782 1993 908
rect 1974 582 1977 588
rect 1978 568 1982 571
rect 1982 542 1985 548
rect 1928 503 1930 507
rect 1934 503 1937 507
rect 1942 503 1944 507
rect 1894 352 1897 368
rect 1942 342 1945 348
rect 1830 322 1833 328
rect 1838 292 1841 318
rect 1928 303 1930 307
rect 1934 303 1937 307
rect 1942 303 1944 307
rect 1990 292 1993 778
rect 2014 752 2017 1148
rect 2022 1132 2025 1158
rect 2030 1042 2033 1078
rect 2054 1062 2057 1328
rect 2062 1282 2065 1378
rect 2102 1362 2105 1378
rect 2070 1352 2073 1358
rect 2126 1312 2129 1878
rect 2150 1772 2153 2158
rect 2158 1982 2161 2068
rect 2166 1952 2169 2928
rect 2174 2912 2177 2998
rect 2182 2622 2185 3098
rect 2250 2788 2257 2791
rect 2222 2692 2225 2738
rect 2230 2662 2233 2738
rect 2174 2002 2177 2438
rect 2186 2348 2190 2351
rect 2182 2302 2185 2308
rect 2198 2162 2201 2248
rect 2166 1932 2169 1948
rect 2162 1798 2166 1801
rect 2138 1638 2145 1641
rect 2142 1572 2145 1638
rect 2150 1562 2153 1748
rect 2022 962 2025 968
rect 2050 958 2054 961
rect 2046 902 2049 948
rect 2030 742 2033 758
rect 2038 752 2041 778
rect 2046 672 2049 748
rect 2010 528 2014 531
rect 2022 522 2025 568
rect 1998 492 2001 518
rect 1998 382 2001 468
rect 2006 372 2009 478
rect 1982 252 1985 268
rect 2006 172 2009 178
rect 1926 158 1934 161
rect 1926 152 1929 158
rect 2014 132 2017 508
rect 2050 478 2054 481
rect 2030 392 2033 448
rect 2026 388 2030 391
rect 2054 362 2057 368
rect 2038 152 2041 218
rect 2046 132 2049 338
rect 1928 103 1930 107
rect 1934 103 1937 107
rect 1942 103 1944 107
rect 1734 72 1737 98
rect 2006 52 2009 98
rect 2046 82 2049 128
rect 2054 72 2057 158
rect 2062 141 2065 938
rect 2086 882 2089 1308
rect 2094 1052 2097 1308
rect 2106 1238 2110 1241
rect 2134 1222 2137 1338
rect 2154 1318 2161 1321
rect 2142 1232 2145 1258
rect 2086 772 2089 838
rect 2074 758 2078 761
rect 2102 572 2105 1188
rect 2118 1151 2121 1188
rect 2118 1148 2126 1151
rect 2122 1078 2126 1081
rect 2110 712 2113 948
rect 2122 928 2126 931
rect 2110 672 2113 678
rect 2110 452 2113 478
rect 2134 422 2137 1118
rect 2142 982 2145 1038
rect 2158 942 2161 1318
rect 2166 1112 2169 1738
rect 2174 1702 2177 1948
rect 2182 1781 2185 1998
rect 2182 1778 2190 1781
rect 2182 1602 2185 1768
rect 2190 1742 2193 1748
rect 2198 1632 2201 2158
rect 2214 2102 2217 2568
rect 2226 2418 2230 2421
rect 2230 2322 2233 2328
rect 2222 2272 2225 2288
rect 2198 1562 2201 1568
rect 2206 1532 2209 1678
rect 2190 1282 2193 1478
rect 2190 1022 2193 1278
rect 2202 1268 2206 1271
rect 2198 1151 2201 1238
rect 2214 1162 2217 2088
rect 2222 1761 2225 1788
rect 2222 1758 2230 1761
rect 2238 1761 2241 2598
rect 2246 1852 2249 2678
rect 2254 2632 2257 2788
rect 2254 2512 2257 2628
rect 2270 2562 2273 2618
rect 2262 2542 2265 2558
rect 2266 2528 2273 2531
rect 2262 2452 2265 2458
rect 2254 2162 2257 2328
rect 2254 2132 2257 2138
rect 2262 2112 2265 2448
rect 2270 2282 2273 2528
rect 2278 2342 2281 3028
rect 2318 2732 2321 2908
rect 2342 2792 2345 2828
rect 2294 2502 2297 2528
rect 2270 1932 2273 2278
rect 2294 2252 2297 2498
rect 2310 2332 2313 2418
rect 2286 2212 2289 2218
rect 2318 2192 2321 2728
rect 2326 2542 2329 2598
rect 2334 2452 2337 2518
rect 2298 2148 2302 2151
rect 2302 2082 2305 2128
rect 2238 1758 2246 1761
rect 2254 1732 2257 1738
rect 2242 1698 2249 1701
rect 2222 1632 2225 1678
rect 2246 1502 2249 1698
rect 2254 1692 2257 1698
rect 2262 1672 2265 1768
rect 2278 1692 2281 1928
rect 2318 1782 2321 2178
rect 2326 2142 2329 2348
rect 2334 2271 2337 2448
rect 2342 2332 2345 2788
rect 2350 2532 2353 2648
rect 2358 2462 2361 2498
rect 2370 2458 2377 2461
rect 2374 2452 2377 2458
rect 2354 2438 2361 2441
rect 2358 2412 2361 2438
rect 2334 2268 2342 2271
rect 2262 1412 2265 1418
rect 2222 1182 2225 1278
rect 2238 1182 2241 1198
rect 2238 1162 2241 1178
rect 2270 1171 2273 1208
rect 2266 1168 2273 1171
rect 2278 1172 2281 1688
rect 2302 1512 2305 1558
rect 2302 1492 2305 1508
rect 2318 1362 2321 1778
rect 2326 1552 2329 2108
rect 2334 2082 2337 2268
rect 2374 2262 2377 2448
rect 2398 2332 2401 2708
rect 2406 2612 2409 3088
rect 2440 3003 2442 3007
rect 2446 3003 2449 3007
rect 2454 3003 2456 3007
rect 2414 2902 2417 2918
rect 2422 2692 2425 2968
rect 2446 2872 2449 2918
rect 2440 2803 2442 2807
rect 2446 2803 2449 2807
rect 2454 2803 2456 2807
rect 2462 2762 2465 2848
rect 2406 2372 2409 2378
rect 2394 2268 2398 2271
rect 2406 2222 2409 2228
rect 2342 2082 2345 2098
rect 2358 1932 2361 2188
rect 2366 1872 2369 2178
rect 2414 2161 2417 2668
rect 2440 2603 2442 2607
rect 2446 2603 2449 2607
rect 2454 2603 2456 2607
rect 2422 2532 2425 2538
rect 2410 2158 2417 2161
rect 2422 2382 2425 2398
rect 2378 2078 2385 2081
rect 2382 1912 2385 2078
rect 2414 2061 2417 2128
rect 2410 2058 2417 2061
rect 2358 1741 2361 1818
rect 2354 1738 2361 1741
rect 2342 1482 2345 1518
rect 2346 1388 2350 1391
rect 2294 1282 2297 1338
rect 2286 1262 2289 1268
rect 2198 1148 2206 1151
rect 2198 1132 2201 1138
rect 2222 1132 2225 1148
rect 2246 1118 2254 1121
rect 2198 1092 2201 1108
rect 2246 1022 2249 1118
rect 2282 1048 2286 1051
rect 2246 962 2249 1018
rect 2222 872 2225 878
rect 2174 742 2177 858
rect 2270 772 2273 1048
rect 2286 822 2289 838
rect 2294 782 2297 1278
rect 2302 812 2305 1288
rect 2318 1222 2321 1358
rect 2330 1348 2334 1351
rect 2350 1172 2353 1348
rect 2358 1082 2361 1738
rect 2366 1722 2369 1868
rect 2406 1802 2409 1818
rect 2366 1542 2369 1718
rect 2378 1648 2382 1651
rect 2382 1492 2385 1618
rect 2422 1602 2425 2378
rect 2430 2342 2433 2408
rect 2440 2403 2442 2407
rect 2446 2403 2449 2407
rect 2454 2403 2456 2407
rect 2462 2342 2465 2358
rect 2470 2312 2473 3018
rect 2478 2512 2481 2518
rect 2486 2462 2489 2638
rect 2494 2432 2497 2608
rect 2502 2562 2505 3098
rect 2502 2552 2505 2558
rect 2482 2358 2486 2361
rect 2440 2203 2442 2207
rect 2446 2203 2449 2207
rect 2454 2203 2456 2207
rect 2442 2068 2446 2071
rect 2440 2003 2442 2007
rect 2446 2003 2449 2007
rect 2454 2003 2456 2007
rect 2430 1902 2433 1928
rect 2478 1872 2481 1878
rect 2440 1803 2442 1807
rect 2446 1803 2449 1807
rect 2454 1803 2456 1807
rect 2462 1802 2465 1848
rect 2458 1758 2462 1761
rect 2440 1603 2442 1607
rect 2446 1603 2449 1607
rect 2454 1603 2456 1607
rect 2470 1542 2473 1858
rect 2462 1538 2470 1541
rect 2422 1512 2425 1528
rect 2382 1392 2385 1488
rect 2402 1468 2406 1471
rect 2390 1112 2393 1458
rect 2414 1452 2417 1468
rect 2406 1282 2409 1318
rect 2414 1292 2417 1448
rect 2440 1403 2442 1407
rect 2446 1403 2449 1407
rect 2454 1403 2456 1407
rect 2398 1092 2401 1128
rect 2318 1052 2321 1078
rect 2358 982 2361 1078
rect 2406 1072 2409 1278
rect 2422 1112 2425 1358
rect 2430 1272 2433 1308
rect 2440 1203 2442 1207
rect 2446 1203 2449 1207
rect 2454 1203 2456 1207
rect 2370 1048 2374 1051
rect 2390 902 2393 908
rect 2314 868 2318 871
rect 2190 722 2193 758
rect 2302 742 2305 808
rect 2350 752 2353 898
rect 2222 738 2230 741
rect 2158 542 2161 718
rect 2190 702 2193 718
rect 2206 642 2209 668
rect 2222 592 2225 738
rect 2358 722 2361 738
rect 2310 672 2313 698
rect 2318 672 2321 688
rect 2230 638 2238 641
rect 2174 572 2177 578
rect 2206 562 2209 568
rect 2102 382 2105 418
rect 2130 388 2137 391
rect 2078 142 2081 148
rect 2062 138 2070 141
rect 2086 92 2089 328
rect 2118 302 2121 328
rect 2134 272 2137 388
rect 2094 132 2097 228
rect 2118 212 2121 218
rect 2118 142 2121 208
rect 2126 82 2129 158
rect 1418 18 1422 21
rect 2090 18 2094 21
rect 2150 11 2153 478
rect 2230 362 2233 638
rect 2238 402 2241 608
rect 2262 492 2265 508
rect 2314 448 2318 451
rect 2342 442 2345 458
rect 2214 122 2217 178
rect 2222 142 2225 148
rect 2238 72 2241 398
rect 2246 342 2249 428
rect 2334 382 2337 438
rect 2262 292 2265 348
rect 2270 282 2273 288
rect 2262 192 2265 198
rect 2286 192 2289 248
rect 2286 32 2289 188
rect 2302 82 2305 368
rect 2326 182 2329 188
rect 2334 112 2337 248
rect 2350 132 2353 488
rect 2374 472 2377 878
rect 2406 872 2409 1028
rect 2430 982 2433 1078
rect 2440 1003 2442 1007
rect 2446 1003 2449 1007
rect 2454 1003 2456 1007
rect 2386 758 2393 761
rect 2358 292 2361 458
rect 2390 442 2393 758
rect 2398 742 2401 768
rect 2406 712 2409 858
rect 2414 802 2417 918
rect 2440 803 2442 807
rect 2446 803 2449 807
rect 2454 803 2456 807
rect 2390 352 2393 438
rect 2398 322 2401 398
rect 2406 372 2409 708
rect 2414 642 2417 648
rect 2422 612 2425 648
rect 2440 603 2442 607
rect 2446 603 2449 607
rect 2454 603 2456 607
rect 2422 592 2425 598
rect 2462 472 2465 1538
rect 2494 1442 2497 2338
rect 2502 2272 2505 2278
rect 2510 2232 2513 2978
rect 2558 2892 2561 2928
rect 2582 2902 2585 2908
rect 2542 2572 2545 2708
rect 2534 2538 2542 2541
rect 2534 2532 2537 2538
rect 2518 1882 2521 2468
rect 2538 2238 2542 2241
rect 2542 2122 2545 2218
rect 2550 2072 2553 2528
rect 2558 2472 2561 2888
rect 2570 2738 2577 2741
rect 2574 2632 2577 2738
rect 2574 2362 2577 2368
rect 2582 2352 2585 2898
rect 2590 2692 2593 2718
rect 2598 2532 2601 2728
rect 2598 2482 2601 2518
rect 2558 2172 2561 2308
rect 2558 2132 2561 2148
rect 2526 2052 2529 2058
rect 2510 1782 2513 1818
rect 2494 1392 2497 1438
rect 2482 1378 2486 1381
rect 2506 1258 2513 1261
rect 2510 1252 2513 1258
rect 2518 1052 2521 1788
rect 2526 1392 2529 1418
rect 2550 1352 2553 1988
rect 2574 1972 2577 2158
rect 2582 2132 2585 2138
rect 2582 1672 2585 2128
rect 2590 1952 2593 2128
rect 2606 1962 2609 3098
rect 2806 2952 2809 2968
rect 2874 2948 2878 2951
rect 2906 2928 2910 2931
rect 2750 2912 2753 2918
rect 2750 2882 2753 2908
rect 2758 2852 2761 2928
rect 2882 2888 2886 2891
rect 2650 2738 2654 2741
rect 2622 2091 2625 2718
rect 2630 2652 2633 2698
rect 2630 2572 2633 2648
rect 2638 2482 2641 2528
rect 2646 2412 2649 2548
rect 2638 2341 2641 2378
rect 2646 2372 2649 2408
rect 2634 2338 2641 2341
rect 2618 2088 2625 2091
rect 2654 2122 2657 2678
rect 2670 2662 2673 2818
rect 2662 2372 2665 2528
rect 2678 2482 2681 2748
rect 2734 2702 2737 2768
rect 2750 2752 2753 2848
rect 2742 2742 2745 2748
rect 2750 2662 2753 2748
rect 2742 2642 2745 2658
rect 2750 2622 2753 2658
rect 2686 2522 2689 2528
rect 2670 2342 2673 2348
rect 2678 2332 2681 2358
rect 2694 2331 2697 2518
rect 2690 2328 2697 2331
rect 2694 2322 2697 2328
rect 2702 2312 2705 2468
rect 2630 2002 2633 2018
rect 2638 2012 2641 2038
rect 2634 1958 2638 1961
rect 2590 1662 2593 1758
rect 2590 1642 2593 1658
rect 2566 1542 2569 1608
rect 2598 1552 2601 1618
rect 2574 1548 2582 1551
rect 2574 1542 2577 1548
rect 2590 1528 2598 1531
rect 2558 1492 2561 1518
rect 2590 1412 2593 1528
rect 2606 1492 2609 1918
rect 2654 1842 2657 2118
rect 2662 1982 2665 2038
rect 2670 1932 2673 2148
rect 2714 2088 2718 2091
rect 2678 2032 2681 2088
rect 2698 2068 2702 2071
rect 2646 1792 2649 1838
rect 2654 1702 2657 1808
rect 2686 1732 2689 2068
rect 2726 1942 2729 2578
rect 2750 2472 2753 2618
rect 2750 2402 2753 2448
rect 2758 2432 2761 2848
rect 2766 2662 2769 2668
rect 2794 2648 2801 2651
rect 2750 2232 2753 2398
rect 2766 2282 2769 2548
rect 2778 2458 2782 2461
rect 2798 2442 2801 2648
rect 2806 2552 2809 2768
rect 2910 2752 2913 2788
rect 2818 2748 2822 2751
rect 2918 2662 2921 2718
rect 2918 2652 2921 2658
rect 2798 2361 2801 2368
rect 2794 2358 2801 2361
rect 2758 2262 2761 2278
rect 2766 2232 2769 2278
rect 2750 2072 2753 2228
rect 2742 2018 2750 2021
rect 2758 2021 2761 2068
rect 2754 2018 2761 2021
rect 2766 2022 2769 2048
rect 2734 2002 2737 2018
rect 2742 1992 2745 2018
rect 2766 1922 2769 2018
rect 2774 1902 2777 2348
rect 2806 2132 2809 2508
rect 2814 2462 2817 2628
rect 2822 2612 2825 2618
rect 2822 2582 2825 2608
rect 2822 2332 2825 2438
rect 2834 2388 2838 2391
rect 2794 2128 2798 2131
rect 2782 2052 2785 2058
rect 2790 1972 2793 2078
rect 2782 1952 2785 1958
rect 2790 1782 2793 1868
rect 2706 1758 2713 1761
rect 2622 1542 2625 1548
rect 2526 1292 2529 1298
rect 2534 1272 2537 1298
rect 2590 1252 2593 1358
rect 2606 1272 2609 1328
rect 2622 1222 2625 1328
rect 2570 1158 2574 1161
rect 2478 492 2481 1048
rect 2510 951 2513 958
rect 2506 948 2513 951
rect 2486 742 2489 858
rect 2502 782 2505 938
rect 2486 598 2494 601
rect 2462 432 2465 468
rect 2486 422 2489 598
rect 2378 268 2382 271
rect 2414 262 2417 348
rect 2422 302 2425 408
rect 2440 403 2442 407
rect 2446 403 2449 407
rect 2454 403 2456 407
rect 2490 388 2494 391
rect 2414 252 2417 258
rect 2358 162 2361 248
rect 2462 212 2465 228
rect 2440 203 2442 207
rect 2446 203 2449 207
rect 2454 203 2456 207
rect 2358 112 2361 158
rect 2426 138 2430 141
rect 2494 132 2497 138
rect 2174 12 2177 28
rect 2502 12 2505 768
rect 2518 751 2521 1048
rect 2526 882 2529 938
rect 2518 748 2526 751
rect 2510 732 2513 738
rect 2522 728 2526 731
rect 2522 718 2526 721
rect 2534 512 2537 1078
rect 2550 1062 2553 1068
rect 2558 982 2561 1148
rect 2590 1082 2593 1188
rect 2598 988 2606 991
rect 2586 878 2590 881
rect 2566 812 2569 828
rect 2598 822 2601 988
rect 2630 962 2633 1368
rect 2638 1312 2641 1328
rect 2638 992 2641 1128
rect 2618 878 2625 881
rect 2622 852 2625 878
rect 2630 862 2633 958
rect 2542 582 2545 808
rect 2550 502 2553 728
rect 2530 448 2534 451
rect 2510 242 2513 448
rect 2518 402 2521 448
rect 2518 352 2521 398
rect 2534 371 2537 378
rect 2530 368 2537 371
rect 2558 292 2561 448
rect 2566 412 2569 748
rect 2598 732 2601 738
rect 2622 692 2625 818
rect 2638 752 2641 988
rect 2622 662 2625 678
rect 2582 552 2585 658
rect 2590 592 2593 658
rect 2610 558 2614 561
rect 2566 348 2574 351
rect 2566 332 2569 348
rect 2566 292 2569 328
rect 2530 178 2534 181
rect 2550 131 2553 228
rect 2546 128 2553 131
rect 2562 128 2566 131
rect 2606 72 2609 88
rect 2630 12 2633 638
rect 2646 392 2649 1678
rect 2654 1662 2657 1698
rect 2686 1242 2689 1728
rect 2710 1702 2713 1758
rect 2750 1692 2753 1738
rect 2738 1688 2742 1691
rect 2766 1691 2769 1758
rect 2766 1688 2774 1691
rect 2710 1648 2718 1651
rect 2710 1242 2713 1648
rect 2718 1462 2721 1548
rect 2726 1462 2729 1468
rect 2742 1292 2745 1408
rect 2734 1272 2737 1278
rect 2654 1122 2657 1128
rect 2738 1118 2742 1121
rect 2702 1092 2705 1118
rect 2766 1112 2769 1688
rect 2790 1592 2793 1638
rect 2786 1528 2790 1531
rect 2778 1268 2782 1271
rect 2790 1152 2793 1358
rect 2798 1331 2801 1998
rect 2806 1932 2809 2128
rect 2814 1962 2817 2318
rect 2842 2218 2846 2221
rect 2878 2192 2881 2408
rect 2834 2148 2838 2151
rect 2826 2138 2830 2141
rect 2862 2092 2865 2108
rect 2886 2092 2889 2588
rect 2830 2081 2833 2088
rect 2826 2078 2833 2081
rect 2814 1882 2817 1908
rect 2822 1562 2825 2038
rect 2902 1752 2905 1938
rect 2926 1882 2929 3008
rect 2952 2903 2954 2907
rect 2958 2903 2961 2907
rect 2966 2903 2968 2907
rect 2934 2562 2937 2738
rect 2942 2672 2945 2728
rect 2952 2703 2954 2707
rect 2958 2703 2961 2707
rect 2966 2703 2968 2707
rect 2974 2602 2977 2958
rect 2990 2722 2993 2728
rect 2998 2702 3001 2738
rect 3006 2672 3009 2808
rect 2942 2512 2945 2538
rect 2974 2532 2977 2598
rect 3006 2562 3009 2668
rect 2952 2503 2954 2507
rect 2958 2503 2961 2507
rect 2966 2503 2968 2507
rect 2974 2362 2977 2528
rect 2998 2472 3001 2478
rect 2952 2303 2954 2307
rect 2958 2303 2961 2307
rect 2966 2303 2968 2307
rect 3006 2262 3009 2548
rect 3014 2302 3017 2378
rect 2994 2168 2998 2171
rect 2952 2103 2954 2107
rect 2958 2103 2961 2107
rect 2966 2103 2968 2107
rect 2942 1942 2945 1948
rect 2952 1903 2954 1907
rect 2958 1903 2961 1907
rect 2966 1903 2968 1907
rect 2974 1882 2977 1898
rect 3010 1838 3014 1841
rect 2952 1703 2954 1707
rect 2958 1703 2961 1707
rect 2966 1703 2968 1707
rect 2830 1632 2833 1648
rect 2870 1642 2873 1648
rect 2822 1542 2825 1558
rect 2830 1522 2833 1628
rect 2878 1602 2881 1638
rect 2798 1328 2809 1331
rect 2798 1282 2801 1318
rect 2678 912 2681 938
rect 2666 878 2670 881
rect 2654 762 2657 848
rect 2662 772 2665 808
rect 2670 802 2673 828
rect 2654 612 2657 758
rect 2678 752 2681 908
rect 2678 592 2681 738
rect 2694 712 2697 728
rect 2654 512 2657 568
rect 2678 561 2681 588
rect 2678 558 2686 561
rect 2654 402 2657 508
rect 2658 178 2665 181
rect 2662 132 2665 178
rect 2670 82 2673 508
rect 2678 482 2681 518
rect 2702 282 2705 1068
rect 2774 1062 2777 1078
rect 2710 562 2713 808
rect 2726 722 2729 758
rect 2722 718 2726 721
rect 2722 658 2726 661
rect 2706 148 2710 151
rect 2694 132 2697 148
rect 2718 82 2721 148
rect 2742 12 2745 978
rect 2750 952 2753 1008
rect 2750 732 2753 948
rect 2774 872 2777 948
rect 2766 842 2769 868
rect 2758 502 2761 728
rect 2766 392 2769 838
rect 2774 772 2777 868
rect 2798 682 2801 868
rect 2806 862 2809 1328
rect 2814 1162 2817 1488
rect 2830 1472 2833 1478
rect 2822 1462 2825 1468
rect 2822 1132 2825 1158
rect 2774 562 2777 598
rect 2774 462 2777 518
rect 2774 452 2777 458
rect 2814 292 2817 1128
rect 2830 1122 2833 1468
rect 2838 1392 2841 1558
rect 2850 1518 2854 1521
rect 2870 1462 2873 1488
rect 2846 1392 2849 1428
rect 2842 1328 2846 1331
rect 2822 561 2825 818
rect 2822 558 2830 561
rect 2830 382 2833 548
rect 2838 302 2841 1208
rect 2854 1172 2857 1418
rect 2862 1052 2865 1108
rect 2854 772 2857 818
rect 2870 532 2873 1298
rect 2878 1152 2881 1578
rect 2886 1551 2889 1598
rect 2886 1548 2894 1551
rect 2898 1458 2902 1461
rect 2886 1432 2889 1438
rect 2902 1272 2905 1458
rect 2902 1172 2905 1218
rect 2878 1012 2881 1148
rect 2886 1082 2889 1088
rect 2886 902 2889 938
rect 2886 852 2889 878
rect 2894 862 2897 978
rect 2902 832 2905 848
rect 2878 712 2881 718
rect 2886 712 2889 798
rect 2894 692 2897 828
rect 2902 632 2905 828
rect 2910 762 2913 1618
rect 2926 1302 2929 1678
rect 2978 1618 2985 1621
rect 2982 1582 2985 1618
rect 2942 1512 2945 1518
rect 2952 1503 2954 1507
rect 2958 1503 2961 1507
rect 2966 1503 2968 1507
rect 2974 1402 2977 1498
rect 2982 1492 2985 1508
rect 2934 1072 2937 1398
rect 2952 1303 2954 1307
rect 2958 1303 2961 1307
rect 2966 1303 2968 1307
rect 2974 1292 2977 1298
rect 2942 1112 2945 1258
rect 2952 1103 2954 1107
rect 2958 1103 2961 1107
rect 2966 1103 2968 1107
rect 2974 1072 2977 1218
rect 2990 1132 2993 1708
rect 3014 1352 3017 1458
rect 3014 1132 3017 1348
rect 3006 1122 3009 1128
rect 2998 1112 3001 1118
rect 2982 1092 2985 1108
rect 2942 1052 2945 1058
rect 2998 1012 3001 1038
rect 3014 1002 3017 1088
rect 3022 1012 3025 3028
rect 3062 2662 3065 2668
rect 3054 2632 3057 2648
rect 3030 2292 3033 2328
rect 3038 2292 3041 2378
rect 3030 1472 3033 2288
rect 3062 2082 3065 2448
rect 3054 1532 3057 1818
rect 3062 1802 3065 2078
rect 3070 1542 3073 2948
rect 3342 2942 3345 2958
rect 3354 2868 3358 2871
rect 3094 2742 3097 2868
rect 3246 2732 3249 2748
rect 3254 2742 3257 2838
rect 3194 2728 3198 2731
rect 3110 2352 3113 2698
rect 3194 2658 3198 2661
rect 3078 2342 3081 2348
rect 3086 2282 3089 2348
rect 3126 2252 3129 2628
rect 3134 2362 3137 2448
rect 3106 2078 3110 2081
rect 3126 2032 3129 2238
rect 3134 2102 3137 2358
rect 3146 2268 3150 2271
rect 3158 2162 3161 2658
rect 3234 2548 3238 2551
rect 3222 2522 3225 2538
rect 3238 2472 3241 2548
rect 3254 2522 3257 2558
rect 3270 2532 3273 2548
rect 3202 2468 3206 2471
rect 3190 2452 3193 2468
rect 3166 2342 3169 2358
rect 3174 2192 3177 2418
rect 3166 2088 3174 2091
rect 3094 1972 3097 2018
rect 3082 1958 3086 1961
rect 3142 1948 3150 1951
rect 3142 1942 3145 1948
rect 3078 1932 3081 1938
rect 3150 1932 3153 1938
rect 3166 1912 3169 2088
rect 3182 1972 3185 2328
rect 3190 2092 3193 2448
rect 3206 2331 3209 2348
rect 3234 2338 3238 2341
rect 3202 2328 3209 2331
rect 3086 1632 3089 1708
rect 3094 1622 3097 1758
rect 3106 1718 3110 1721
rect 3030 1372 3033 1468
rect 3094 1402 3097 1618
rect 3102 1562 3105 1618
rect 3118 1512 3121 1748
rect 3182 1742 3185 1938
rect 3130 1728 3134 1731
rect 3154 1658 3161 1661
rect 3158 1652 3161 1658
rect 3166 1652 3169 1678
rect 3182 1632 3185 1648
rect 3126 1592 3129 1618
rect 3110 1452 3113 1468
rect 3066 1288 3073 1291
rect 3046 1162 3049 1278
rect 3070 1232 3073 1288
rect 3062 1192 3065 1198
rect 3058 1158 3062 1161
rect 2918 822 2921 918
rect 2952 903 2954 907
rect 2958 903 2961 907
rect 2966 903 2968 907
rect 2942 872 2945 898
rect 2934 852 2937 858
rect 2918 762 2921 818
rect 2894 592 2897 628
rect 2918 622 2921 668
rect 2926 652 2929 848
rect 2974 822 2977 838
rect 2952 703 2954 707
rect 2958 703 2961 707
rect 2966 703 2968 707
rect 2952 503 2954 507
rect 2958 503 2961 507
rect 2966 503 2968 507
rect 2954 488 2958 491
rect 2974 472 2977 708
rect 2990 662 2993 698
rect 3006 652 3009 658
rect 2926 442 2929 448
rect 2894 352 2897 358
rect 2806 272 2809 278
rect 2806 102 2809 268
rect 2862 252 2865 338
rect 2926 302 2929 328
rect 2934 272 2937 298
rect 2858 248 2862 251
rect 2942 212 2945 308
rect 2952 303 2954 307
rect 2958 303 2961 307
rect 2966 303 2968 307
rect 2974 212 2977 468
rect 2990 362 2993 648
rect 2998 512 3001 628
rect 3006 452 3009 648
rect 3022 452 3025 848
rect 3054 352 3057 458
rect 3062 392 3065 1018
rect 3070 942 3073 1148
rect 3078 1131 3081 1178
rect 3102 1152 3105 1158
rect 3110 1148 3118 1151
rect 3110 1142 3113 1148
rect 3078 1128 3086 1131
rect 3090 1078 3094 1081
rect 3110 1072 3113 1078
rect 3086 912 3089 1038
rect 3086 892 3089 908
rect 3118 902 3121 948
rect 3126 912 3129 978
rect 3134 962 3137 1608
rect 3166 1572 3169 1578
rect 3190 1532 3193 1798
rect 3198 1532 3201 2228
rect 3230 2152 3233 2208
rect 3238 2182 3241 2208
rect 3206 2032 3209 2148
rect 3214 2142 3217 2148
rect 3246 2092 3249 2458
rect 3254 2372 3257 2518
rect 3278 2482 3281 2528
rect 3270 2192 3273 2438
rect 3254 2082 3257 2088
rect 3238 2052 3241 2078
rect 3214 1952 3217 1958
rect 3222 1902 3225 1998
rect 3258 1938 3262 1941
rect 3278 1932 3281 2478
rect 3362 2468 3369 2471
rect 3326 2462 3329 2468
rect 3310 2412 3313 2458
rect 3302 2252 3305 2268
rect 3286 2151 3289 2178
rect 3286 2148 3294 2151
rect 3310 2112 3313 2408
rect 3298 2048 3302 2051
rect 3318 1942 3321 2458
rect 3366 2422 3369 2468
rect 3350 2262 3353 2278
rect 3338 2258 3342 2261
rect 3334 2052 3337 2068
rect 3350 2052 3353 2258
rect 3358 2152 3361 2338
rect 3382 2271 3385 3048
rect 3472 3003 3474 3007
rect 3478 3003 3481 3007
rect 3486 3003 3488 3007
rect 3402 2928 3406 2931
rect 3390 2922 3393 2928
rect 3490 2888 3497 2891
rect 3494 2872 3497 2888
rect 3472 2803 3474 2807
rect 3478 2803 3481 2807
rect 3486 2803 3488 2807
rect 3474 2768 3478 2771
rect 3390 2532 3393 2548
rect 3422 2532 3425 2728
rect 3430 2682 3433 2748
rect 3502 2742 3505 2988
rect 3526 2862 3529 3018
rect 3942 2962 3945 3038
rect 3710 2942 3713 2948
rect 3542 2752 3545 2908
rect 3550 2832 3553 2878
rect 3574 2822 3577 2878
rect 3506 2738 3510 2741
rect 3472 2603 3474 2607
rect 3478 2603 3481 2607
rect 3486 2603 3488 2607
rect 3582 2562 3585 2888
rect 3590 2842 3593 2868
rect 3382 2268 3393 2271
rect 3370 2258 3374 2261
rect 3342 1952 3345 1968
rect 3346 1948 3350 1951
rect 3214 1662 3217 1758
rect 3278 1732 3281 1928
rect 3246 1642 3249 1648
rect 3206 1552 3209 1558
rect 3146 1528 3150 1531
rect 3170 1528 3174 1531
rect 3182 1528 3190 1531
rect 3166 1282 3169 1518
rect 3174 1282 3177 1338
rect 3150 1161 3153 1258
rect 3166 1172 3169 1278
rect 3182 1272 3185 1528
rect 3198 1222 3201 1368
rect 3214 1362 3217 1628
rect 3222 1472 3225 1478
rect 3222 1272 3225 1288
rect 3206 1162 3209 1178
rect 3150 1158 3158 1161
rect 3142 1082 3145 1148
rect 3150 1122 3153 1128
rect 3134 952 3137 958
rect 3150 942 3153 988
rect 3098 888 3102 891
rect 3118 891 3121 898
rect 3118 888 3126 891
rect 3158 862 3161 1148
rect 3198 1022 3201 1128
rect 3070 672 3073 838
rect 3078 812 3081 828
rect 3110 732 3113 738
rect 3054 242 3057 288
rect 2952 103 2954 107
rect 2958 103 2961 107
rect 2966 103 2968 107
rect 2974 82 2977 88
rect 3078 82 3081 628
rect 3118 562 3121 778
rect 3094 462 3097 478
rect 3118 472 3121 478
rect 3094 442 3097 448
rect 3102 252 3105 278
rect 3118 182 3121 438
rect 3134 292 3137 788
rect 3158 712 3161 858
rect 3158 482 3161 588
rect 3166 561 3169 828
rect 3174 722 3177 888
rect 3182 842 3185 868
rect 3190 842 3193 858
rect 3198 832 3201 838
rect 3206 802 3209 1078
rect 3166 558 3174 561
rect 3198 522 3201 638
rect 3214 592 3217 1228
rect 3238 1222 3241 1538
rect 3270 1362 3273 1658
rect 3278 1482 3281 1728
rect 3294 1572 3297 1758
rect 3302 1652 3305 1698
rect 3310 1562 3313 1588
rect 3334 1562 3337 1898
rect 3318 1532 3321 1558
rect 3314 1478 3318 1481
rect 3278 1352 3281 1478
rect 3298 1468 3302 1471
rect 3326 1471 3329 1548
rect 3350 1532 3353 1538
rect 3338 1528 3342 1531
rect 3366 1531 3369 1548
rect 3362 1528 3369 1531
rect 3374 1522 3377 1528
rect 3326 1468 3334 1471
rect 3334 1452 3337 1468
rect 3358 1452 3361 1478
rect 3370 1468 3377 1471
rect 3374 1452 3377 1468
rect 3382 1462 3385 1968
rect 3390 1702 3393 2268
rect 3398 2262 3401 2278
rect 3406 2062 3409 2418
rect 3422 2292 3425 2528
rect 3502 2442 3505 2518
rect 3534 2462 3537 2478
rect 3542 2462 3545 2478
rect 3522 2458 3526 2461
rect 3472 2403 3474 2407
rect 3478 2403 3481 2407
rect 3486 2403 3488 2407
rect 3406 1822 3409 2058
rect 3414 2052 3417 2068
rect 3422 1782 3425 2248
rect 3430 2202 3433 2288
rect 3472 2203 3474 2207
rect 3478 2203 3481 2207
rect 3486 2203 3488 2207
rect 3494 2202 3497 2428
rect 3554 2338 3561 2341
rect 3570 2338 3577 2341
rect 3542 2268 3550 2271
rect 3542 2152 3545 2268
rect 3558 2212 3561 2338
rect 3574 2242 3577 2338
rect 3514 2068 3518 2071
rect 3462 2012 3465 2048
rect 3472 2003 3474 2007
rect 3478 2003 3481 2007
rect 3486 2003 3488 2007
rect 3414 1712 3417 1748
rect 3322 1448 3326 1451
rect 3250 1338 3257 1341
rect 3254 1272 3257 1338
rect 3254 1262 3257 1268
rect 3226 1128 3230 1131
rect 3238 1042 3241 1208
rect 3246 1122 3249 1238
rect 3254 1142 3257 1148
rect 3278 1082 3281 1348
rect 3306 1338 3313 1341
rect 3286 1322 3289 1328
rect 3310 1312 3313 1338
rect 3354 1338 3358 1341
rect 3342 1332 3345 1338
rect 3330 1328 3337 1331
rect 3302 1172 3305 1198
rect 3238 862 3241 988
rect 3246 872 3249 1058
rect 3262 902 3265 1058
rect 3230 848 3238 851
rect 3286 851 3289 1078
rect 3318 962 3321 1328
rect 3298 928 3302 931
rect 3310 922 3313 928
rect 3318 902 3321 958
rect 3278 848 3289 851
rect 3230 682 3233 848
rect 3246 672 3249 708
rect 3262 692 3265 698
rect 3262 652 3265 688
rect 3238 592 3241 608
rect 3214 541 3217 558
rect 3210 538 3217 541
rect 3166 462 3169 488
rect 3142 232 3145 288
rect 3174 282 3177 478
rect 3182 472 3185 488
rect 3214 412 3217 538
rect 3250 528 3254 531
rect 3230 462 3233 508
rect 3230 362 3233 378
rect 3254 341 3257 358
rect 3262 352 3265 398
rect 3278 392 3281 848
rect 3286 652 3289 838
rect 3298 788 3302 791
rect 3302 692 3305 738
rect 3302 592 3305 688
rect 3326 572 3329 1308
rect 3334 1052 3337 1328
rect 3366 1242 3369 1268
rect 3334 862 3337 1048
rect 3342 562 3345 1008
rect 3350 922 3353 938
rect 3358 702 3361 1048
rect 3366 692 3369 768
rect 3374 672 3377 1418
rect 3390 1392 3393 1698
rect 3422 1662 3425 1778
rect 3430 1722 3433 1998
rect 3434 1718 3441 1721
rect 3398 1552 3401 1558
rect 3414 1522 3417 1548
rect 3398 1252 3401 1278
rect 3406 1262 3409 1468
rect 3414 1442 3417 1518
rect 3426 1468 3430 1471
rect 3438 1422 3441 1718
rect 3446 1682 3449 1718
rect 3454 1692 3457 1908
rect 3494 1882 3497 1898
rect 3472 1803 3474 1807
rect 3478 1803 3481 1807
rect 3486 1803 3488 1807
rect 3510 1702 3513 1938
rect 3526 1902 3529 2108
rect 3542 1932 3545 2148
rect 3518 1852 3521 1888
rect 3526 1872 3529 1888
rect 3526 1772 3529 1808
rect 3426 1298 3430 1301
rect 3422 1288 3430 1291
rect 3390 1122 3393 1238
rect 3398 951 3401 1138
rect 3422 1112 3425 1288
rect 3434 1268 3438 1271
rect 3446 1192 3449 1208
rect 3454 1181 3457 1688
rect 3482 1678 3486 1681
rect 3470 1642 3473 1648
rect 3502 1642 3505 1688
rect 3472 1603 3474 1607
rect 3478 1603 3481 1607
rect 3486 1603 3488 1607
rect 3462 1512 3465 1578
rect 3502 1532 3505 1538
rect 3510 1532 3513 1698
rect 3574 1552 3577 2078
rect 3590 2002 3593 2688
rect 3598 2552 3601 2898
rect 3638 2832 3641 2878
rect 3614 2682 3617 2828
rect 3630 2732 3633 2788
rect 3654 2721 3657 2818
rect 3654 2718 3662 2721
rect 3654 2692 3657 2718
rect 3606 2582 3609 2588
rect 3598 2512 3601 2548
rect 3622 2492 3625 2518
rect 3670 2462 3673 2878
rect 3694 2732 3697 2928
rect 3690 2598 3697 2601
rect 3694 2572 3697 2598
rect 3658 2428 3662 2431
rect 3606 2242 3609 2418
rect 3614 2072 3617 2378
rect 3598 1802 3601 1928
rect 3546 1548 3550 1551
rect 3582 1542 3585 1558
rect 3590 1532 3593 1728
rect 3530 1528 3534 1531
rect 3474 1508 3478 1511
rect 3472 1403 3474 1407
rect 3478 1403 3481 1407
rect 3486 1403 3488 1407
rect 3472 1203 3474 1207
rect 3478 1203 3481 1207
rect 3486 1203 3488 1207
rect 3454 1178 3462 1181
rect 3482 1148 3486 1151
rect 3494 1151 3497 1398
rect 3502 1312 3505 1518
rect 3546 1488 3550 1491
rect 3526 1212 3529 1368
rect 3542 1352 3545 1358
rect 3558 1332 3561 1518
rect 3598 1432 3601 1648
rect 3606 1352 3609 1958
rect 3614 1942 3617 2068
rect 3646 1982 3649 2068
rect 3614 1742 3617 1938
rect 3614 1512 3617 1738
rect 3622 1682 3625 1858
rect 3654 1852 3657 2238
rect 3654 1762 3657 1848
rect 3630 1541 3633 1758
rect 3670 1752 3673 2458
rect 3686 2272 3689 2328
rect 3642 1658 3649 1661
rect 3626 1538 3633 1541
rect 3622 1422 3625 1528
rect 3610 1348 3617 1351
rect 3542 1152 3545 1328
rect 3598 1272 3601 1338
rect 3558 1172 3561 1178
rect 3494 1148 3502 1151
rect 3502 1132 3505 1148
rect 3450 1078 3454 1081
rect 3470 1052 3473 1058
rect 3526 1042 3529 1118
rect 3472 1003 3474 1007
rect 3478 1003 3481 1007
rect 3486 1003 3488 1007
rect 3394 948 3401 951
rect 3414 932 3417 938
rect 3422 922 3425 928
rect 3402 858 3406 861
rect 3362 658 3366 661
rect 3294 512 3297 528
rect 3350 492 3353 628
rect 3310 462 3313 468
rect 3326 392 3329 408
rect 3382 352 3385 748
rect 3422 701 3425 708
rect 3418 698 3425 701
rect 3434 698 3438 701
rect 3390 661 3393 688
rect 3390 658 3398 661
rect 3250 338 3257 341
rect 2974 72 2977 78
rect 3174 72 3177 258
rect 3246 192 3249 338
rect 3406 302 3409 608
rect 3414 531 3417 688
rect 3454 662 3457 968
rect 3498 838 3505 841
rect 3502 822 3505 838
rect 3472 803 3474 807
rect 3478 803 3481 807
rect 3486 803 3488 807
rect 3414 528 3422 531
rect 3406 292 3409 298
rect 3422 232 3425 528
rect 3454 292 3457 658
rect 3462 552 3465 758
rect 3502 742 3505 818
rect 3514 718 3518 721
rect 3502 642 3505 678
rect 3472 603 3474 607
rect 3478 603 3481 607
rect 3486 603 3488 607
rect 3518 552 3521 568
rect 3462 352 3465 548
rect 3472 403 3474 407
rect 3478 403 3481 407
rect 3486 403 3488 407
rect 3494 362 3497 408
rect 3470 242 3473 248
rect 3358 162 3361 198
rect 3422 172 3425 228
rect 3454 192 3457 238
rect 3518 222 3521 328
rect 3526 322 3529 898
rect 3542 892 3545 1088
rect 3566 1062 3569 1178
rect 3574 1082 3577 1198
rect 3582 1192 3585 1238
rect 3574 1032 3577 1068
rect 3594 1058 3598 1061
rect 3590 922 3593 928
rect 3542 672 3545 728
rect 3550 482 3553 888
rect 3566 792 3569 808
rect 3566 772 3569 788
rect 3598 622 3601 1038
rect 3606 782 3609 1198
rect 3614 1142 3617 1348
rect 3622 1282 3625 1318
rect 3622 1262 3625 1278
rect 3630 1191 3633 1438
rect 3626 1188 3633 1191
rect 3606 762 3609 778
rect 3614 762 3617 1138
rect 3622 1092 3625 1188
rect 3622 1012 3625 1088
rect 3622 962 3625 1008
rect 3630 992 3633 1148
rect 3622 772 3625 938
rect 3614 652 3617 758
rect 3630 692 3633 988
rect 3638 751 3641 1548
rect 3646 1442 3649 1658
rect 3646 1342 3649 1348
rect 3646 1042 3649 1248
rect 3654 951 3657 1748
rect 3678 1712 3681 1958
rect 3694 1832 3697 2468
rect 3702 2302 3705 2718
rect 3718 2562 3721 2888
rect 3726 2882 3729 2918
rect 3726 2732 3729 2878
rect 3742 2752 3745 2958
rect 3718 2542 3721 2558
rect 3726 2432 3729 2728
rect 3758 2722 3761 2738
rect 3742 2642 3745 2658
rect 3758 2542 3761 2718
rect 3766 2562 3769 2928
rect 3798 2772 3801 2788
rect 3710 2132 3713 2138
rect 3710 2052 3713 2088
rect 3718 1952 3721 2148
rect 3734 2142 3737 2388
rect 3742 2232 3745 2268
rect 3774 2182 3777 2618
rect 3790 2512 3793 2768
rect 3830 2541 3833 2738
rect 3838 2728 3846 2731
rect 3838 2722 3841 2728
rect 3830 2538 3838 2541
rect 3834 2528 3838 2531
rect 3790 2412 3793 2508
rect 3846 2502 3849 2628
rect 3854 2522 3857 2578
rect 3818 2338 3822 2341
rect 3862 2332 3865 2858
rect 3918 2822 3921 2868
rect 3870 2332 3873 2338
rect 3894 2332 3897 2528
rect 3910 2482 3913 2778
rect 3902 2352 3905 2358
rect 3854 2282 3857 2298
rect 3778 2148 3782 2151
rect 3798 2042 3801 2158
rect 3822 2082 3825 2088
rect 3846 2062 3849 2208
rect 3862 2192 3865 2328
rect 3886 2072 3889 2298
rect 3918 2282 3921 2288
rect 3934 2232 3937 2908
rect 3942 2842 3945 2958
rect 3976 2903 3978 2907
rect 3982 2903 3985 2907
rect 3990 2903 3992 2907
rect 4030 2852 4033 3048
rect 4098 2988 4105 2991
rect 4102 2752 4105 2988
rect 3958 2732 3961 2748
rect 4062 2742 4065 2748
rect 3966 2682 3969 2718
rect 3998 2712 4001 2728
rect 4094 2722 4097 2728
rect 3976 2703 3978 2707
rect 3982 2703 3985 2707
rect 3990 2703 3992 2707
rect 3998 2622 4001 2698
rect 4086 2692 4089 2718
rect 4038 2632 4041 2668
rect 3966 2372 3969 2508
rect 3976 2503 3978 2507
rect 3982 2503 3985 2507
rect 3990 2503 3992 2507
rect 3976 2303 3978 2307
rect 3982 2303 3985 2307
rect 3990 2303 3992 2307
rect 4006 2282 4009 2568
rect 4022 2362 4025 2608
rect 4038 2582 4041 2628
rect 4086 2622 4089 2688
rect 4102 2652 4105 2748
rect 4110 2732 4113 3028
rect 4130 2958 4134 2961
rect 4142 2792 4145 2998
rect 4150 2952 4153 2958
rect 4122 2738 4126 2741
rect 4134 2652 4137 2758
rect 4134 2572 4137 2648
rect 3986 2278 3990 2281
rect 3958 2072 3961 2108
rect 3810 2058 3814 2061
rect 3894 2061 3897 2068
rect 3890 2058 3897 2061
rect 3710 1862 3713 1888
rect 3702 1792 3705 1828
rect 3694 1651 3697 1668
rect 3690 1648 3697 1651
rect 3702 1572 3705 1728
rect 3690 1528 3694 1531
rect 3710 1492 3713 1818
rect 3666 1338 3670 1341
rect 3678 1282 3681 1478
rect 3690 1278 3694 1281
rect 3718 1252 3721 1948
rect 3726 1742 3729 1868
rect 3734 1862 3737 1888
rect 3742 1792 3745 1938
rect 3750 1892 3753 1918
rect 3754 1858 3758 1861
rect 3734 1492 3737 1778
rect 3742 1512 3745 1788
rect 3750 1772 3753 1818
rect 3766 1751 3769 1968
rect 3798 1882 3801 1928
rect 3766 1748 3774 1751
rect 3762 1738 3766 1741
rect 3750 1672 3753 1678
rect 3762 1538 3769 1541
rect 3766 1532 3769 1538
rect 3694 1162 3697 1198
rect 3710 1162 3713 1178
rect 3726 1152 3729 1218
rect 3678 1062 3681 1138
rect 3654 948 3662 951
rect 3662 771 3665 878
rect 3658 768 3665 771
rect 3638 748 3646 751
rect 3638 732 3641 738
rect 3686 692 3689 858
rect 3566 582 3569 598
rect 3598 482 3601 608
rect 3598 281 3601 468
rect 3614 352 3617 588
rect 3694 492 3697 1118
rect 3710 1062 3713 1088
rect 3718 1002 3721 1108
rect 3742 1082 3745 1358
rect 3750 1172 3753 1288
rect 3758 1262 3761 1438
rect 3782 1362 3785 1768
rect 3790 1712 3793 1758
rect 3774 1262 3777 1268
rect 3782 1172 3785 1328
rect 3798 1322 3801 1868
rect 3806 1472 3809 2058
rect 3846 1932 3849 2058
rect 3902 1908 3910 1911
rect 3814 1591 3817 1878
rect 3826 1848 3830 1851
rect 3830 1691 3833 1698
rect 3826 1688 3833 1691
rect 3814 1588 3822 1591
rect 3834 1558 3838 1561
rect 3834 1548 3838 1551
rect 3758 1132 3761 1138
rect 3702 862 3705 878
rect 3710 862 3713 968
rect 3718 892 3721 968
rect 3726 772 3729 1078
rect 3738 1068 3742 1071
rect 3754 938 3758 941
rect 3766 932 3769 948
rect 3774 942 3777 1168
rect 3782 1152 3785 1168
rect 3710 692 3713 728
rect 3702 662 3705 668
rect 3718 591 3721 748
rect 3774 652 3777 938
rect 3782 662 3785 798
rect 3718 588 3726 591
rect 3726 512 3729 588
rect 3774 542 3777 648
rect 3790 582 3793 1068
rect 3806 832 3809 1468
rect 3830 1052 3833 1478
rect 3870 1252 3873 1288
rect 3878 1282 3881 1908
rect 3886 1572 3889 1888
rect 3902 1712 3905 1908
rect 3910 1442 3913 1888
rect 3918 1762 3921 1838
rect 3926 1622 3929 1678
rect 3926 1542 3929 1618
rect 3934 1562 3937 1578
rect 3942 1482 3945 2008
rect 3950 1962 3953 2068
rect 3950 1652 3953 1678
rect 3910 1262 3913 1438
rect 3818 1028 3822 1031
rect 3818 938 3822 941
rect 3806 742 3809 758
rect 3726 462 3729 508
rect 3674 438 3678 441
rect 3698 358 3702 361
rect 3686 302 3689 318
rect 3594 278 3601 281
rect 3472 203 3474 207
rect 3478 203 3481 207
rect 3486 203 3488 207
rect 3458 168 3462 171
rect 3182 122 3185 128
rect 3350 92 3353 118
rect 3174 62 3177 68
rect 3374 52 3377 98
rect 3574 91 3577 178
rect 3570 88 3577 91
rect 3590 92 3593 258
rect 3638 182 3641 248
rect 3654 132 3657 278
rect 3710 222 3713 378
rect 3722 338 3726 341
rect 3718 211 3721 218
rect 3714 208 3721 211
rect 3726 212 3729 318
rect 3742 292 3745 398
rect 3798 372 3801 588
rect 3750 342 3753 348
rect 3734 131 3737 208
rect 3814 152 3817 488
rect 3822 462 3825 758
rect 3830 742 3833 1048
rect 3838 822 3841 1008
rect 3862 892 3865 1198
rect 3882 1128 3886 1131
rect 3942 1082 3945 1478
rect 3950 1452 3953 1568
rect 3958 1112 3961 1198
rect 3958 1062 3961 1068
rect 3846 752 3849 868
rect 3898 858 3905 861
rect 3902 842 3905 858
rect 3822 352 3825 458
rect 3826 228 3833 231
rect 3830 212 3833 228
rect 3830 152 3833 208
rect 3838 142 3841 418
rect 3854 372 3857 378
rect 3862 142 3865 728
rect 3870 542 3873 698
rect 3878 672 3881 678
rect 3894 572 3897 838
rect 3902 702 3905 838
rect 3910 742 3913 918
rect 3958 892 3961 958
rect 3926 852 3929 868
rect 3934 752 3937 758
rect 3902 582 3905 648
rect 3902 522 3905 558
rect 3934 542 3937 548
rect 3894 402 3897 448
rect 3886 332 3889 378
rect 3886 222 3889 308
rect 3894 262 3897 398
rect 3910 342 3913 358
rect 3902 231 3905 238
rect 3898 228 3905 231
rect 3734 128 3742 131
rect 3798 102 3801 128
rect 3590 72 3593 88
rect 3726 72 3729 88
rect 3806 82 3809 118
rect 3902 82 3905 198
rect 3918 192 3921 528
rect 3938 368 3942 371
rect 3926 282 3929 348
rect 3958 342 3961 608
rect 3966 332 3969 2138
rect 3976 2103 3978 2107
rect 3982 2103 3985 2107
rect 3990 2103 3992 2107
rect 3998 1952 4001 2148
rect 3976 1903 3978 1907
rect 3982 1903 3985 1907
rect 3990 1903 3992 1907
rect 3976 1703 3978 1707
rect 3982 1703 3985 1707
rect 3990 1703 3992 1707
rect 3976 1503 3978 1507
rect 3982 1503 3985 1507
rect 3990 1503 3992 1507
rect 3998 1442 4001 1948
rect 4006 1852 4009 2068
rect 4014 2032 4017 2218
rect 4022 2072 4025 2188
rect 4030 2092 4033 2328
rect 4030 2042 4033 2068
rect 4038 1952 4041 2318
rect 4054 2152 4057 2488
rect 4134 2482 4137 2568
rect 4142 2552 4145 2788
rect 4150 2542 4153 2648
rect 4062 2302 4065 2378
rect 4062 2172 4065 2248
rect 4046 2072 4049 2078
rect 4038 1802 4041 1818
rect 4046 1772 4049 2038
rect 4046 1732 4049 1768
rect 4054 1752 4057 2148
rect 4062 2102 4065 2168
rect 4074 2158 4078 2161
rect 4078 2102 4081 2128
rect 4062 2082 4065 2088
rect 4074 2068 4078 2071
rect 4062 1912 4065 2048
rect 4030 1652 4033 1728
rect 4046 1652 4049 1728
rect 4046 1522 4049 1558
rect 4014 1362 4017 1378
rect 4050 1368 4054 1371
rect 3976 1303 3978 1307
rect 3982 1303 3985 1307
rect 3990 1303 3992 1307
rect 3998 1152 4001 1158
rect 3976 1103 3978 1107
rect 3982 1103 3985 1107
rect 3990 1103 3992 1107
rect 3998 912 4001 928
rect 3976 903 3978 907
rect 3982 903 3985 907
rect 3990 903 3992 907
rect 4006 732 4009 918
rect 3976 703 3978 707
rect 3982 703 3985 707
rect 3990 703 3992 707
rect 3976 503 3978 507
rect 3982 503 3985 507
rect 3990 503 3992 507
rect 4006 482 4009 728
rect 4002 468 4006 471
rect 3958 312 3961 328
rect 3974 322 3977 328
rect 3976 303 3978 307
rect 3982 303 3985 307
rect 3990 303 3992 307
rect 3966 282 3969 298
rect 3926 142 3929 268
rect 3976 103 3978 107
rect 3982 103 3985 107
rect 3990 103 3992 107
rect 3682 68 3686 71
rect 3726 62 3729 68
rect 3998 62 4001 418
rect 4014 252 4017 1268
rect 4022 1052 4025 1258
rect 4022 552 4025 668
rect 4030 332 4033 348
rect 4038 112 4041 1368
rect 4050 1248 4054 1251
rect 4062 1242 4065 1908
rect 4054 1152 4057 1178
rect 4054 802 4057 968
rect 4046 768 4054 771
rect 4046 642 4049 768
rect 4062 762 4065 1058
rect 4070 1012 4073 1118
rect 4054 502 4057 748
rect 4062 642 4065 748
rect 4078 672 4081 1938
rect 4086 1772 4089 2128
rect 4094 1952 4097 2288
rect 4150 2262 4153 2268
rect 4102 2142 4105 2148
rect 4114 2078 4118 2081
rect 4134 1968 4142 1971
rect 4110 1861 4113 1868
rect 4106 1858 4113 1861
rect 4086 1382 4089 1458
rect 4086 992 4089 1118
rect 4078 572 4081 648
rect 4074 558 4078 561
rect 4086 462 4089 568
rect 4078 392 4081 448
rect 4062 222 4065 358
rect 4070 262 4073 308
rect 4082 268 4086 271
rect 4070 172 4073 228
rect 4094 112 4097 1438
rect 4102 1032 4105 1738
rect 4110 1672 4113 1758
rect 4122 1648 4126 1651
rect 4134 1641 4137 1968
rect 4142 1882 4145 1888
rect 4150 1802 4153 2028
rect 4142 1652 4145 1688
rect 4134 1638 4145 1641
rect 4122 1358 4126 1361
rect 4118 1348 4126 1351
rect 4134 1351 4137 1478
rect 4130 1348 4137 1351
rect 4118 1282 4121 1348
rect 4142 1232 4145 1638
rect 4150 1332 4153 1348
rect 4158 1262 4161 3058
rect 4166 2492 4169 3068
rect 4174 2802 4177 3048
rect 4174 2472 4177 2708
rect 4166 2102 4169 2288
rect 4174 2081 4177 2458
rect 4170 2078 4177 2081
rect 4166 1882 4169 1968
rect 4174 1932 4177 1938
rect 4170 1758 4174 1761
rect 4170 1538 4174 1541
rect 4182 1372 4185 3038
rect 4190 2942 4193 2958
rect 4190 2872 4193 2938
rect 4190 2632 4193 2868
rect 4190 1572 4193 2488
rect 4198 1732 4201 3078
rect 4250 3068 4254 3071
rect 4230 3062 4233 3068
rect 4266 3048 4270 3051
rect 4278 3042 4281 3068
rect 4302 3032 4305 3048
rect 4218 2948 4222 2951
rect 4206 2672 4209 2708
rect 4206 2342 4209 2608
rect 4214 2452 4217 2928
rect 4246 2772 4249 2998
rect 4238 2752 4241 2758
rect 4242 2738 4246 2741
rect 4214 2281 4217 2388
rect 4210 2278 4217 2281
rect 4222 2132 4225 2578
rect 4190 1422 4193 1558
rect 4198 1482 4201 1728
rect 4110 882 4113 948
rect 4118 792 4121 938
rect 4126 802 4129 868
rect 4106 758 4110 761
rect 4118 752 4121 788
rect 4110 532 4113 558
rect 4102 122 4105 428
rect 4118 232 4121 448
rect 4134 62 4137 1068
rect 4146 1058 4150 1061
rect 4158 1061 4161 1158
rect 4158 1058 4166 1061
rect 4150 852 4153 878
rect 4142 152 4145 558
rect 4150 432 4153 828
rect 4158 102 4161 1048
rect 4166 822 4169 1048
rect 4174 1032 4177 1328
rect 4182 952 4185 1348
rect 4190 1082 4193 1418
rect 4198 1072 4201 1188
rect 4198 962 4201 1068
rect 4174 402 4177 558
rect 4174 272 4177 278
rect 4150 92 4153 98
rect 4142 82 4145 88
rect 4174 52 4177 108
rect 4182 72 4185 948
rect 4190 862 4193 888
rect 4198 882 4201 958
rect 4206 882 4209 1948
rect 4222 1902 4225 2078
rect 4214 1292 4217 1478
rect 4222 1292 4225 1898
rect 4230 1702 4233 2708
rect 4238 2032 4241 2478
rect 4254 2312 4257 2928
rect 4262 2432 4265 3018
rect 4262 2282 4265 2408
rect 4270 2352 4273 2848
rect 4238 1852 4241 2008
rect 4254 1942 4257 1958
rect 4230 1462 4233 1468
rect 4238 1462 4241 1848
rect 4250 1748 4254 1751
rect 4246 1682 4249 1708
rect 4214 1271 4217 1288
rect 4214 1268 4222 1271
rect 4222 1092 4225 1158
rect 4222 1022 4225 1028
rect 4214 962 4217 968
rect 4198 762 4201 878
rect 4206 782 4209 868
rect 4190 462 4193 568
rect 4198 212 4201 758
rect 4214 442 4217 658
rect 4206 192 4209 358
rect 4222 262 4225 1008
rect 4230 712 4233 1318
rect 4238 1072 4241 1238
rect 4246 1052 4249 1548
rect 4254 1352 4257 1748
rect 4262 1672 4265 1928
rect 4266 1468 4270 1471
rect 4242 1038 4246 1041
rect 4246 952 4249 958
rect 4254 942 4257 1328
rect 4270 1042 4273 1118
rect 4246 742 4249 858
rect 4230 441 4233 568
rect 4230 438 4238 441
rect 4238 292 4241 358
rect 4254 292 4257 778
rect 4262 552 4265 938
rect 4270 912 4273 1018
rect 4270 552 4273 748
rect 4278 662 4281 2738
rect 4286 1802 4289 2768
rect 4294 2752 4297 2758
rect 4294 2532 4297 2648
rect 4294 2262 4297 2268
rect 4294 1892 4297 1968
rect 4286 1592 4289 1648
rect 4294 1362 4297 1778
rect 4302 1732 4305 2998
rect 4318 2731 4321 3088
rect 4334 2752 4337 2968
rect 4330 2738 4334 2741
rect 4318 2728 4329 2731
rect 4310 2562 4313 2718
rect 4310 2542 4313 2558
rect 4318 2352 4321 2688
rect 4302 1622 4305 1718
rect 4310 1632 4313 1958
rect 4310 1471 4313 1608
rect 4306 1468 4313 1471
rect 4286 1202 4289 1238
rect 4286 1162 4289 1168
rect 4294 1152 4297 1358
rect 4294 1052 4297 1148
rect 4302 1132 4305 1458
rect 4310 1092 4313 1338
rect 4286 862 4289 938
rect 4270 532 4273 548
rect 4262 232 4265 388
rect 4278 352 4281 658
rect 4286 542 4289 848
rect 4286 352 4289 358
rect 4294 182 4297 1048
rect 4310 852 4313 868
rect 4302 642 4305 648
rect 4302 262 4305 428
rect 4298 158 4302 161
rect 4298 148 4302 151
rect 4302 132 4305 138
rect 4202 88 4206 91
rect 4310 62 4313 668
rect 4318 142 4321 2338
rect 4326 2132 4329 2728
rect 4326 2072 4329 2098
rect 4326 1592 4329 1868
rect 4334 1832 4337 2078
rect 4342 1952 4345 2648
rect 4350 2322 4353 3058
rect 4358 2372 4361 2798
rect 4366 2452 4369 3018
rect 4374 2562 4377 2698
rect 4342 1922 4345 1948
rect 4326 1062 4329 1568
rect 4334 1272 4337 1798
rect 4342 1792 4345 1918
rect 4334 861 4337 1118
rect 4342 1082 4345 1778
rect 4350 1112 4353 2308
rect 4366 2152 4369 2428
rect 4382 2372 4385 2688
rect 4358 1782 4361 2098
rect 4366 2082 4369 2148
rect 4374 2102 4377 2358
rect 4382 2091 4385 2348
rect 4374 2088 4385 2091
rect 4358 1632 4361 1698
rect 4366 1652 4369 2058
rect 4366 1112 4369 1638
rect 4334 858 4345 861
rect 4334 562 4337 848
rect 4342 572 4345 858
rect 4358 672 4361 1088
rect 4330 448 4334 451
rect 4342 182 4345 478
rect 4358 382 4361 668
rect 4366 612 4369 848
rect 4374 312 4377 2088
rect 4390 1752 4393 2688
rect 4386 1308 4393 1311
rect 4390 1082 4393 1308
rect 4362 158 4366 161
rect 4322 128 4326 131
rect 4382 82 4385 748
rect 4322 68 4326 71
rect 4170 38 4174 41
rect 2150 8 2158 11
rect 392 3 394 7
rect 398 3 401 7
rect 406 3 408 7
rect 1416 3 1418 7
rect 1422 3 1425 7
rect 1430 3 1432 7
rect 2440 3 2442 7
rect 2446 3 2449 7
rect 2454 3 2456 7
rect 3472 3 3474 7
rect 3478 3 3481 7
rect 3486 3 3488 7
<< m5contact >>
rect 898 3103 902 3107
rect 905 3103 906 3107
rect 906 3103 909 3107
rect 1930 3103 1934 3107
rect 1937 3103 1938 3107
rect 1938 3103 1941 3107
rect 2954 3103 2958 3107
rect 2961 3103 2962 3107
rect 2962 3103 2965 3107
rect 3978 3103 3982 3107
rect 3985 3103 3986 3107
rect 3986 3103 3989 3107
rect 222 3068 226 3072
rect 630 3068 634 3072
rect 318 3058 322 3062
rect 394 3003 398 3007
rect 401 3003 402 3007
rect 402 3003 405 3007
rect 30 2148 34 2152
rect 14 1788 18 1792
rect 118 2558 122 2562
rect 182 2168 186 2172
rect 190 2148 194 2152
rect 158 1938 162 1942
rect 166 1738 170 1742
rect 158 1678 162 1682
rect 182 1938 186 1942
rect 702 3058 706 3062
rect 394 2803 398 2807
rect 401 2803 402 2807
rect 402 2803 405 2807
rect 394 2603 398 2607
rect 401 2603 402 2607
rect 402 2603 405 2607
rect 394 2403 398 2407
rect 401 2403 402 2407
rect 402 2403 405 2407
rect 394 2203 398 2207
rect 401 2203 402 2207
rect 402 2203 405 2207
rect 366 2038 370 2042
rect 394 2003 398 2007
rect 401 2003 402 2007
rect 402 2003 405 2007
rect 190 1928 194 1932
rect 294 1888 298 1892
rect 390 1868 394 1872
rect 394 1803 398 1807
rect 401 1803 402 1807
rect 402 1803 405 1807
rect 394 1603 398 1607
rect 401 1603 402 1607
rect 402 1603 405 1607
rect 78 1438 82 1442
rect 22 1278 26 1282
rect 14 1238 18 1242
rect 22 1178 26 1182
rect 174 1468 178 1472
rect 430 1918 434 1922
rect 198 1458 202 1462
rect 394 1403 398 1407
rect 401 1403 402 1407
rect 402 1403 405 1407
rect 110 1348 114 1352
rect 246 1328 250 1332
rect 394 1203 398 1207
rect 401 1203 402 1207
rect 402 1203 405 1207
rect 134 688 138 692
rect 166 1068 170 1072
rect 166 868 170 872
rect 166 738 170 742
rect 214 338 218 342
rect 214 148 218 152
rect 394 1003 398 1007
rect 401 1003 402 1007
rect 402 1003 405 1007
rect 158 88 162 92
rect 394 803 398 807
rect 401 803 402 807
rect 402 803 405 807
rect 390 668 394 672
rect 394 603 398 607
rect 401 603 402 607
rect 402 603 405 607
rect 526 2048 530 2052
rect 534 1878 538 1882
rect 550 1678 554 1682
rect 510 1468 514 1472
rect 510 1318 514 1322
rect 502 1258 506 1262
rect 526 1338 530 1342
rect 534 1258 538 1262
rect 574 2558 578 2562
rect 590 1798 594 1802
rect 606 1718 610 1722
rect 518 968 522 972
rect 394 403 398 407
rect 401 403 402 407
rect 402 403 405 407
rect 646 2088 650 2092
rect 646 2058 650 2062
rect 590 1518 594 1522
rect 598 1478 602 1482
rect 606 1458 610 1462
rect 646 1468 650 1472
rect 898 2903 902 2907
rect 905 2903 906 2907
rect 906 2903 909 2907
rect 798 2748 802 2752
rect 1006 2748 1010 2752
rect 898 2703 902 2707
rect 905 2703 906 2707
rect 906 2703 909 2707
rect 830 2528 834 2532
rect 822 2458 826 2462
rect 814 2258 818 2262
rect 806 2158 810 2162
rect 814 2138 818 2142
rect 702 2048 706 2052
rect 726 1968 730 1972
rect 718 1938 722 1942
rect 678 1898 682 1902
rect 726 1858 730 1862
rect 718 1778 722 1782
rect 718 1688 722 1692
rect 710 1438 714 1442
rect 774 2048 778 2052
rect 758 1468 762 1472
rect 766 1358 770 1362
rect 670 1288 674 1292
rect 678 1278 682 1282
rect 694 1188 698 1192
rect 686 1158 690 1162
rect 654 1128 658 1132
rect 662 958 666 962
rect 750 1328 754 1332
rect 702 1068 706 1072
rect 758 1178 762 1182
rect 750 1148 754 1152
rect 798 1808 802 1812
rect 898 2503 902 2507
rect 905 2503 906 2507
rect 906 2503 909 2507
rect 898 2303 902 2307
rect 905 2303 906 2307
rect 906 2303 909 2307
rect 838 2258 842 2262
rect 822 1888 826 1892
rect 822 1768 826 1772
rect 790 1648 794 1652
rect 814 1628 818 1632
rect 814 1548 818 1552
rect 838 2158 842 2162
rect 846 2148 850 2152
rect 838 1888 842 1892
rect 846 1878 850 1882
rect 854 1788 858 1792
rect 870 1908 874 1912
rect 870 1878 874 1882
rect 918 2148 922 2152
rect 1038 2258 1042 2262
rect 902 2138 906 2142
rect 898 2103 902 2107
rect 905 2103 906 2107
rect 906 2103 909 2107
rect 918 1938 922 1942
rect 898 1903 902 1907
rect 905 1903 906 1907
rect 906 1903 909 1907
rect 910 1828 914 1832
rect 910 1728 914 1732
rect 898 1703 902 1707
rect 905 1703 906 1707
rect 906 1703 909 1707
rect 1014 2138 1018 2142
rect 998 1968 1002 1972
rect 998 1858 1002 1862
rect 1022 1978 1026 1982
rect 838 1478 842 1482
rect 894 1548 898 1552
rect 878 1528 882 1532
rect 838 1378 842 1382
rect 806 1208 810 1212
rect 774 1048 778 1052
rect 758 858 762 862
rect 898 1503 902 1507
rect 905 1503 906 1507
rect 906 1503 909 1507
rect 886 1488 890 1492
rect 918 1358 922 1362
rect 926 1338 930 1342
rect 918 1318 922 1322
rect 898 1303 902 1307
rect 905 1303 906 1307
rect 906 1303 909 1307
rect 926 1268 930 1272
rect 926 1238 930 1242
rect 926 1198 930 1202
rect 926 1158 930 1162
rect 974 1688 978 1692
rect 966 1348 970 1352
rect 982 1568 986 1572
rect 934 1148 938 1152
rect 814 868 818 872
rect 822 848 826 852
rect 898 1103 902 1107
rect 905 1103 906 1107
rect 906 1103 909 1107
rect 934 1078 938 1082
rect 898 903 902 907
rect 905 903 906 907
rect 906 903 909 907
rect 534 278 538 282
rect 394 203 398 207
rect 401 203 402 207
rect 402 203 405 207
rect 494 168 498 172
rect 550 58 554 62
rect 774 398 778 402
rect 898 703 902 707
rect 905 703 906 707
rect 906 703 909 707
rect 918 688 922 692
rect 942 668 946 672
rect 1030 1468 1034 1472
rect 1086 2318 1090 2322
rect 1070 2058 1074 2062
rect 1078 1648 1082 1652
rect 1118 2338 1122 2342
rect 1142 1978 1146 1982
rect 1134 1958 1138 1962
rect 1142 1928 1146 1932
rect 1134 1898 1138 1902
rect 1118 1888 1122 1892
rect 1134 1868 1138 1872
rect 1134 1798 1138 1802
rect 1174 2048 1178 2052
rect 1174 1968 1178 1972
rect 1142 1718 1146 1722
rect 1134 1668 1138 1672
rect 1166 1668 1170 1672
rect 1118 1648 1122 1652
rect 1006 1318 1010 1322
rect 974 1128 978 1132
rect 982 1068 986 1072
rect 974 848 978 852
rect 726 318 730 322
rect 898 503 902 507
rect 905 503 906 507
rect 906 503 909 507
rect 1054 1238 1058 1242
rect 1046 1088 1050 1092
rect 1038 1018 1042 1022
rect 1022 898 1026 902
rect 1038 978 1042 982
rect 1094 1508 1098 1512
rect 1102 1478 1106 1482
rect 1102 1288 1106 1292
rect 1078 1208 1082 1212
rect 1070 1158 1074 1162
rect 1078 1068 1082 1072
rect 1102 1178 1106 1182
rect 1126 1548 1130 1552
rect 1118 1188 1122 1192
rect 1238 1938 1242 1942
rect 1230 1738 1234 1742
rect 1286 2628 1290 2632
rect 1278 1938 1282 1942
rect 1286 1878 1290 1882
rect 1418 3003 1422 3007
rect 1425 3003 1426 3007
rect 1426 3003 1429 3007
rect 1462 2948 1466 2952
rect 1598 2888 1602 2892
rect 1558 2868 1562 2872
rect 1418 2803 1422 2807
rect 1425 2803 1426 2807
rect 1426 2803 1429 2807
rect 1374 2458 1378 2462
rect 1358 2448 1362 2452
rect 1334 2268 1338 2272
rect 1326 2078 1330 2082
rect 1318 2028 1322 2032
rect 1238 1718 1242 1722
rect 1150 1048 1154 1052
rect 1182 1178 1186 1182
rect 1134 948 1138 952
rect 1150 948 1154 952
rect 1142 878 1146 882
rect 1134 738 1138 742
rect 898 303 902 307
rect 905 303 906 307
rect 906 303 909 307
rect 950 298 954 302
rect 918 268 922 272
rect 838 228 842 232
rect 694 158 698 162
rect 990 148 994 152
rect 898 103 902 107
rect 905 103 906 107
rect 906 103 909 107
rect 1286 1768 1290 1772
rect 1302 1728 1306 1732
rect 1278 1688 1282 1692
rect 1214 1358 1218 1362
rect 1206 1298 1210 1302
rect 1198 1148 1202 1152
rect 1206 1138 1210 1142
rect 1206 1108 1210 1112
rect 1206 948 1210 952
rect 1230 1328 1234 1332
rect 1230 1168 1234 1172
rect 1238 1128 1242 1132
rect 1222 958 1226 962
rect 1230 938 1234 942
rect 1198 428 1202 432
rect 1150 318 1154 322
rect 1222 488 1226 492
rect 1278 1348 1282 1352
rect 1262 1338 1266 1342
rect 1326 1908 1330 1912
rect 1318 1808 1322 1812
rect 1350 2098 1354 2102
rect 1334 1618 1338 1622
rect 1326 1368 1330 1372
rect 1342 1378 1346 1382
rect 1418 2603 1422 2607
rect 1425 2603 1426 2607
rect 1426 2603 1429 2607
rect 1510 2538 1514 2542
rect 1446 2448 1450 2452
rect 1518 2408 1522 2412
rect 1418 2403 1422 2407
rect 1425 2403 1426 2407
rect 1426 2403 1429 2407
rect 1398 2348 1402 2352
rect 1366 1968 1370 1972
rect 1374 1848 1378 1852
rect 1382 1748 1386 1752
rect 1382 1718 1386 1722
rect 1382 1688 1386 1692
rect 1366 1658 1370 1662
rect 1366 1568 1370 1572
rect 1374 1538 1378 1542
rect 1350 1338 1354 1342
rect 1310 1318 1314 1322
rect 1342 1308 1346 1312
rect 1294 1258 1298 1262
rect 1326 1248 1330 1252
rect 1278 1128 1282 1132
rect 1270 1098 1274 1102
rect 1262 1078 1266 1082
rect 1254 968 1258 972
rect 1262 948 1266 952
rect 1302 1058 1306 1062
rect 1310 1058 1314 1062
rect 1278 858 1282 862
rect 1358 1218 1362 1222
rect 1350 1078 1354 1082
rect 1334 928 1338 932
rect 1374 1348 1378 1352
rect 1390 1318 1394 1322
rect 1382 1288 1386 1292
rect 1374 1278 1378 1282
rect 1382 1278 1386 1282
rect 1382 1198 1386 1202
rect 1390 1188 1394 1192
rect 1374 1148 1378 1152
rect 1326 918 1330 922
rect 1350 838 1354 842
rect 1310 678 1314 682
rect 1254 668 1258 672
rect 1230 398 1234 402
rect 1198 268 1202 272
rect 1118 158 1122 162
rect 1150 148 1154 152
rect 1118 138 1122 142
rect 1086 128 1090 132
rect 1102 78 1106 82
rect 1214 168 1218 172
rect 1270 298 1274 302
rect 1254 148 1258 152
rect 1278 158 1282 162
rect 1262 128 1266 132
rect 1294 478 1298 482
rect 1310 348 1314 352
rect 1294 338 1298 342
rect 1366 748 1370 752
rect 1350 318 1354 322
rect 1310 188 1314 192
rect 1310 138 1314 142
rect 1254 78 1258 82
rect 1418 2203 1422 2207
rect 1425 2203 1426 2207
rect 1426 2203 1429 2207
rect 1526 2158 1530 2162
rect 1418 2003 1422 2007
rect 1425 2003 1426 2007
rect 1426 2003 1429 2007
rect 1462 1978 1466 1982
rect 1414 1928 1418 1932
rect 1418 1803 1422 1807
rect 1425 1803 1426 1807
rect 1426 1803 1429 1807
rect 1446 1918 1450 1922
rect 1462 1888 1466 1892
rect 1454 1828 1458 1832
rect 1446 1668 1450 1672
rect 1418 1603 1422 1607
rect 1425 1603 1426 1607
rect 1426 1603 1429 1607
rect 1462 1558 1466 1562
rect 1398 1128 1402 1132
rect 1418 1403 1422 1407
rect 1425 1403 1426 1407
rect 1426 1403 1429 1407
rect 1414 1348 1418 1352
rect 1414 1258 1418 1262
rect 1438 1208 1442 1212
rect 1418 1203 1422 1207
rect 1425 1203 1426 1207
rect 1426 1203 1429 1207
rect 1418 1003 1422 1007
rect 1425 1003 1426 1007
rect 1426 1003 1429 1007
rect 1398 898 1402 902
rect 1398 888 1402 892
rect 1398 868 1402 872
rect 1382 818 1386 822
rect 1418 803 1422 807
rect 1425 803 1426 807
rect 1426 803 1429 807
rect 1430 778 1434 782
rect 1422 768 1426 772
rect 1406 648 1410 652
rect 1418 603 1422 607
rect 1425 603 1426 607
rect 1426 603 1429 607
rect 1478 1548 1482 1552
rect 1462 1358 1466 1362
rect 1502 1918 1506 1922
rect 1510 1868 1514 1872
rect 1510 1748 1514 1752
rect 1510 1648 1514 1652
rect 1510 1548 1514 1552
rect 1494 1478 1498 1482
rect 1502 1458 1506 1462
rect 1494 1388 1498 1392
rect 1486 1368 1490 1372
rect 1542 1768 1546 1772
rect 1526 1708 1530 1712
rect 1518 1518 1522 1522
rect 1678 2948 1682 2952
rect 1750 2878 1754 2882
rect 1678 2478 1682 2482
rect 1622 2318 1626 2322
rect 1606 2268 1610 2272
rect 1654 2428 1658 2432
rect 1646 2388 1650 2392
rect 1582 2038 1586 2042
rect 1582 1948 1586 1952
rect 1574 1898 1578 1902
rect 1558 1818 1562 1822
rect 1574 1718 1578 1722
rect 1606 1668 1610 1672
rect 1550 1628 1554 1632
rect 1550 1528 1554 1532
rect 1606 1528 1610 1532
rect 1510 1338 1514 1342
rect 1470 1258 1474 1262
rect 1486 1328 1490 1332
rect 1494 1228 1498 1232
rect 1478 1078 1482 1082
rect 1470 1048 1474 1052
rect 1462 1028 1466 1032
rect 1454 868 1458 872
rect 1454 848 1458 852
rect 1342 88 1346 92
rect 1238 68 1242 72
rect 1334 28 1338 32
rect 1374 128 1378 132
rect 1390 118 1394 122
rect 1414 548 1418 552
rect 1446 478 1450 482
rect 1462 708 1466 712
rect 1462 698 1466 702
rect 1462 558 1466 562
rect 1418 403 1422 407
rect 1425 403 1426 407
rect 1426 403 1429 407
rect 1486 988 1490 992
rect 1526 1378 1530 1382
rect 1558 1498 1562 1502
rect 1550 1338 1554 1342
rect 1526 1318 1530 1322
rect 1550 1308 1554 1312
rect 1542 1298 1546 1302
rect 1542 1248 1546 1252
rect 1534 1228 1538 1232
rect 1566 1418 1570 1422
rect 1574 1348 1578 1352
rect 1590 1448 1594 1452
rect 1638 2048 1642 2052
rect 1678 2458 1682 2462
rect 1702 2438 1706 2442
rect 1702 2278 1706 2282
rect 1662 1868 1666 1872
rect 1670 1868 1674 1872
rect 1694 2088 1698 2092
rect 1670 1758 1674 1762
rect 1646 1608 1650 1612
rect 1638 1568 1642 1572
rect 1750 2588 1754 2592
rect 1734 2478 1738 2482
rect 1718 2258 1722 2262
rect 1726 2058 1730 2062
rect 1758 2358 1762 2362
rect 1814 2548 1818 2552
rect 1806 2528 1810 2532
rect 1806 2488 1810 2492
rect 1766 2348 1770 2352
rect 1782 2348 1786 2352
rect 1758 2178 1762 2182
rect 1750 1968 1754 1972
rect 1750 1958 1754 1962
rect 1766 2168 1770 2172
rect 1766 1888 1770 1892
rect 1718 1878 1722 1882
rect 1718 1868 1722 1872
rect 1742 1858 1746 1862
rect 1758 1858 1762 1862
rect 1718 1738 1722 1742
rect 1678 1648 1682 1652
rect 1654 1558 1658 1562
rect 1678 1518 1682 1522
rect 1614 1358 1618 1362
rect 1598 1348 1602 1352
rect 1574 1328 1578 1332
rect 1574 1178 1578 1182
rect 1558 1128 1562 1132
rect 1534 1118 1538 1122
rect 1534 1088 1538 1092
rect 1542 1078 1546 1082
rect 1510 988 1514 992
rect 1518 988 1522 992
rect 1510 968 1514 972
rect 1566 1088 1570 1092
rect 1590 1278 1594 1282
rect 1614 1318 1618 1322
rect 1686 1478 1690 1482
rect 1638 1448 1642 1452
rect 1646 1408 1650 1412
rect 1654 1408 1658 1412
rect 1638 1358 1642 1362
rect 1638 1308 1642 1312
rect 1606 1278 1610 1282
rect 1622 1278 1626 1282
rect 1550 918 1554 922
rect 1542 908 1546 912
rect 1558 908 1562 912
rect 1494 808 1498 812
rect 1486 658 1490 662
rect 1438 268 1442 272
rect 1550 788 1554 792
rect 1486 388 1490 392
rect 1518 358 1522 362
rect 1486 258 1490 262
rect 1478 238 1482 242
rect 1510 228 1514 232
rect 1418 203 1422 207
rect 1425 203 1426 207
rect 1426 203 1429 207
rect 1406 138 1410 142
rect 1582 838 1586 842
rect 1590 798 1594 802
rect 1582 708 1586 712
rect 1558 618 1562 622
rect 1542 428 1546 432
rect 1630 1178 1634 1182
rect 1622 1128 1626 1132
rect 1622 1108 1626 1112
rect 1622 1068 1626 1072
rect 1678 1438 1682 1442
rect 1670 1348 1674 1352
rect 1662 1088 1666 1092
rect 1654 1038 1658 1042
rect 1638 1028 1642 1032
rect 1654 928 1658 932
rect 1654 868 1658 872
rect 1686 978 1690 982
rect 1686 878 1690 882
rect 1670 828 1674 832
rect 1614 728 1618 732
rect 1614 678 1618 682
rect 1598 598 1602 602
rect 1798 2228 1802 2232
rect 1806 2148 1810 2152
rect 1806 1908 1810 1912
rect 1798 1718 1802 1722
rect 1790 1708 1794 1712
rect 1798 1688 1802 1692
rect 1742 1558 1746 1562
rect 1758 1528 1762 1532
rect 1806 1668 1810 1672
rect 1806 1628 1810 1632
rect 1726 1468 1730 1472
rect 1758 1468 1762 1472
rect 1798 1448 1802 1452
rect 1758 1428 1762 1432
rect 1726 1398 1730 1402
rect 1718 1328 1722 1332
rect 1734 1328 1738 1332
rect 1734 1318 1738 1322
rect 1718 1308 1722 1312
rect 1742 1278 1746 1282
rect 1766 1328 1770 1332
rect 1750 1248 1754 1252
rect 1758 1248 1762 1252
rect 1766 1228 1770 1232
rect 1750 1218 1754 1222
rect 1702 1118 1706 1122
rect 1702 1068 1706 1072
rect 1710 1058 1714 1062
rect 1710 1008 1714 1012
rect 1750 958 1754 962
rect 1798 1258 1802 1262
rect 1782 1218 1786 1222
rect 1774 1098 1778 1102
rect 1774 1088 1778 1092
rect 1766 1068 1770 1072
rect 1726 888 1730 892
rect 1726 878 1730 882
rect 1726 868 1730 872
rect 1702 798 1706 802
rect 1702 738 1706 742
rect 1662 728 1666 732
rect 1694 718 1698 722
rect 1646 708 1650 712
rect 1550 138 1554 142
rect 1438 78 1442 82
rect 1502 78 1506 82
rect 1590 88 1594 92
rect 1382 58 1386 62
rect 1566 58 1570 62
rect 1606 198 1610 202
rect 1606 148 1610 152
rect 1638 138 1642 142
rect 1662 578 1666 582
rect 1718 758 1722 762
rect 1830 2368 1834 2372
rect 1862 2528 1866 2532
rect 1854 2458 1858 2462
rect 1846 2428 1850 2432
rect 1846 2338 1850 2342
rect 1862 2318 1866 2322
rect 1854 2288 1858 2292
rect 1846 2258 1850 2262
rect 1838 2088 1842 2092
rect 1814 1558 1818 1562
rect 1830 2008 1834 2012
rect 1862 2248 1866 2252
rect 1870 2038 1874 2042
rect 1838 1838 1842 1842
rect 1822 1398 1826 1402
rect 1822 1308 1826 1312
rect 1822 1228 1826 1232
rect 1822 1188 1826 1192
rect 1822 1088 1826 1092
rect 1798 788 1802 792
rect 1838 1428 1842 1432
rect 1830 878 1834 882
rect 1930 2903 1934 2907
rect 1937 2903 1938 2907
rect 1938 2903 1941 2907
rect 1930 2703 1934 2707
rect 1937 2703 1938 2707
rect 1938 2703 1941 2707
rect 1894 2638 1898 2642
rect 1930 2503 1934 2507
rect 1937 2503 1938 2507
rect 1938 2503 1941 2507
rect 1950 2498 1954 2502
rect 1918 2478 1922 2482
rect 1910 2448 1914 2452
rect 1886 2018 1890 2022
rect 1930 2303 1934 2307
rect 1937 2303 1938 2307
rect 1938 2303 1941 2307
rect 1930 2103 1934 2107
rect 1937 2103 1938 2107
rect 1938 2103 1941 2107
rect 1982 2908 1986 2912
rect 1982 2658 1986 2662
rect 1966 2288 1970 2292
rect 2046 2618 2050 2622
rect 2014 2568 2018 2572
rect 1982 2358 1986 2362
rect 1998 2338 2002 2342
rect 2054 2438 2058 2442
rect 2062 2358 2066 2362
rect 2014 2298 2018 2302
rect 2014 2278 2018 2282
rect 1990 2248 1994 2252
rect 2006 2248 2010 2252
rect 2022 2248 2026 2252
rect 1982 2228 1986 2232
rect 2006 2178 2010 2182
rect 1998 2138 2002 2142
rect 1950 2038 1954 2042
rect 1966 2018 1970 2022
rect 1950 1988 1954 1992
rect 1934 1968 1938 1972
rect 1910 1938 1914 1942
rect 2054 2168 2058 2172
rect 2062 2028 2066 2032
rect 2094 2688 2098 2692
rect 2094 2648 2098 2652
rect 2086 2578 2090 2582
rect 2086 2528 2090 2532
rect 2086 2458 2090 2462
rect 2158 2878 2162 2882
rect 2078 2368 2082 2372
rect 2094 2348 2098 2352
rect 2110 2298 2114 2302
rect 2142 2408 2146 2412
rect 2126 2258 2130 2262
rect 1934 1928 1938 1932
rect 1894 1858 1898 1862
rect 1878 1778 1882 1782
rect 1886 1718 1890 1722
rect 1870 1618 1874 1622
rect 1886 1578 1890 1582
rect 1870 1568 1874 1572
rect 1886 1518 1890 1522
rect 1894 1498 1898 1502
rect 1894 1478 1898 1482
rect 1870 1368 1874 1372
rect 1878 1358 1882 1362
rect 1886 1278 1890 1282
rect 1854 1078 1858 1082
rect 1862 1078 1866 1082
rect 1854 1058 1858 1062
rect 1854 968 1858 972
rect 1894 1268 1898 1272
rect 1870 918 1874 922
rect 1870 888 1874 892
rect 1854 818 1858 822
rect 1862 808 1866 812
rect 1870 808 1874 812
rect 1774 688 1778 692
rect 1758 468 1762 472
rect 1742 398 1746 402
rect 1678 348 1682 352
rect 1726 348 1730 352
rect 1710 138 1714 142
rect 1774 458 1778 462
rect 1846 698 1850 702
rect 1886 918 1890 922
rect 1854 568 1858 572
rect 1798 368 1802 372
rect 1782 278 1786 282
rect 1930 1903 1934 1907
rect 1937 1903 1938 1907
rect 1938 1903 1941 1907
rect 1990 1778 1994 1782
rect 2014 1738 2018 1742
rect 1974 1728 1978 1732
rect 1958 1708 1962 1712
rect 1930 1703 1934 1707
rect 1937 1703 1938 1707
rect 1938 1703 1941 1707
rect 1926 1668 1930 1672
rect 1918 1638 1922 1642
rect 1974 1628 1978 1632
rect 1910 1478 1914 1482
rect 1910 1428 1914 1432
rect 1966 1598 1970 1602
rect 1966 1588 1970 1592
rect 1926 1528 1930 1532
rect 1930 1503 1934 1507
rect 1937 1503 1938 1507
rect 1938 1503 1941 1507
rect 1926 1438 1930 1442
rect 1926 1418 1930 1422
rect 1942 1378 1946 1382
rect 1910 1308 1914 1312
rect 1930 1303 1934 1307
rect 1937 1303 1938 1307
rect 1938 1303 1941 1307
rect 1902 838 1906 842
rect 1918 1178 1922 1182
rect 1930 1103 1934 1107
rect 1937 1103 1938 1107
rect 1938 1103 1941 1107
rect 1974 1558 1978 1562
rect 1910 808 1914 812
rect 1902 708 1906 712
rect 1902 628 1906 632
rect 1930 903 1934 907
rect 1937 903 1938 907
rect 1938 903 1941 907
rect 1942 848 1946 852
rect 1930 703 1934 707
rect 1937 703 1938 707
rect 1938 703 1941 707
rect 2006 1668 2010 1672
rect 2014 1668 2018 1672
rect 2054 1888 2058 1892
rect 2062 1858 2066 1862
rect 2054 1798 2058 1802
rect 2062 1758 2066 1762
rect 2046 1748 2050 1752
rect 2046 1738 2050 1742
rect 2062 1738 2066 1742
rect 2006 1638 2010 1642
rect 2102 1858 2106 1862
rect 2086 1768 2090 1772
rect 2078 1608 2082 1612
rect 2006 1558 2010 1562
rect 2102 1718 2106 1722
rect 2142 1978 2146 1982
rect 2142 1958 2146 1962
rect 2102 1538 2106 1542
rect 2014 1448 2018 1452
rect 1982 1238 1986 1242
rect 1998 1388 2002 1392
rect 2062 1378 2066 1382
rect 2110 1378 2114 1382
rect 2006 1348 2010 1352
rect 2014 1308 2018 1312
rect 2038 1278 2042 1282
rect 1998 1218 2002 1222
rect 1998 1128 2002 1132
rect 1990 968 1994 972
rect 1974 838 1978 842
rect 1990 778 1994 782
rect 1974 578 1978 582
rect 1982 568 1986 572
rect 1982 548 1986 552
rect 1930 503 1934 507
rect 1937 503 1938 507
rect 1938 503 1941 507
rect 1942 348 1946 352
rect 1830 328 1834 332
rect 1930 303 1934 307
rect 1937 303 1938 307
rect 1938 303 1941 307
rect 2022 1128 2026 1132
rect 2102 1358 2106 1362
rect 2070 1348 2074 1352
rect 2158 1978 2162 1982
rect 2222 2738 2226 2742
rect 2174 2438 2178 2442
rect 2182 2348 2186 2352
rect 2182 2308 2186 2312
rect 2166 1948 2170 1952
rect 2158 1798 2162 1802
rect 2142 1568 2146 1572
rect 2134 1338 2138 1342
rect 2126 1308 2130 1312
rect 2030 1038 2034 1042
rect 2022 968 2026 972
rect 2054 958 2058 962
rect 2046 948 2050 952
rect 2038 748 2042 752
rect 2030 738 2034 742
rect 2014 528 2018 532
rect 1998 518 2002 522
rect 1982 248 1986 252
rect 2006 168 2010 172
rect 1926 148 1930 152
rect 2046 478 2050 482
rect 2022 388 2026 392
rect 2054 368 2058 372
rect 1930 103 1934 107
rect 1937 103 1938 107
rect 1938 103 1941 107
rect 2102 1238 2106 1242
rect 2142 1258 2146 1262
rect 2118 1188 2122 1192
rect 2086 768 2090 772
rect 2070 758 2074 762
rect 2126 1078 2130 1082
rect 2118 928 2122 932
rect 2110 678 2114 682
rect 2110 478 2114 482
rect 2142 1038 2146 1042
rect 2190 1748 2194 1752
rect 2222 2418 2226 2422
rect 2230 2318 2234 2322
rect 2222 2288 2226 2292
rect 2214 2088 2218 2092
rect 2206 1678 2210 1682
rect 2198 1568 2202 1572
rect 2198 1268 2202 1272
rect 2198 1238 2202 1242
rect 2222 1788 2226 1792
rect 2262 2558 2266 2562
rect 2262 2458 2266 2462
rect 2254 2158 2258 2162
rect 2254 2128 2258 2132
rect 2318 2728 2322 2732
rect 2294 2498 2298 2502
rect 2310 2328 2314 2332
rect 2294 2248 2298 2252
rect 2286 2218 2290 2222
rect 2326 2348 2330 2352
rect 2294 2148 2298 2152
rect 2302 2128 2306 2132
rect 2262 1768 2266 1772
rect 2254 1728 2258 1732
rect 2222 1678 2226 1682
rect 2254 1698 2258 1702
rect 2358 2498 2362 2502
rect 2374 2448 2378 2452
rect 2358 2408 2362 2412
rect 2262 1418 2266 1422
rect 2270 1208 2274 1212
rect 2238 1198 2242 1202
rect 2222 1178 2226 1182
rect 2238 1178 2242 1182
rect 2302 1488 2306 1492
rect 2442 3003 2446 3007
rect 2449 3003 2450 3007
rect 2450 3003 2453 3007
rect 2414 2918 2418 2922
rect 2446 2868 2450 2872
rect 2442 2803 2446 2807
rect 2449 2803 2450 2807
rect 2450 2803 2453 2807
rect 2406 2368 2410 2372
rect 2390 2268 2394 2272
rect 2406 2228 2410 2232
rect 2342 2078 2346 2082
rect 2442 2603 2446 2607
rect 2449 2603 2450 2607
rect 2450 2603 2453 2607
rect 2422 2538 2426 2542
rect 2422 2378 2426 2382
rect 2358 1818 2362 1822
rect 2326 1548 2330 1552
rect 2342 1478 2346 1482
rect 2342 1388 2346 1392
rect 2302 1288 2306 1292
rect 2286 1258 2290 1262
rect 2198 1138 2202 1142
rect 2198 1088 2202 1092
rect 2270 1048 2274 1052
rect 2278 1048 2282 1052
rect 2190 1018 2194 1022
rect 2246 958 2250 962
rect 2222 878 2226 882
rect 2174 858 2178 862
rect 2286 838 2290 842
rect 2326 1348 2330 1352
rect 2318 1218 2322 1222
rect 2350 1168 2354 1172
rect 2406 1818 2410 1822
rect 2382 1648 2386 1652
rect 2382 1618 2386 1622
rect 2442 2403 2446 2407
rect 2449 2403 2450 2407
rect 2450 2403 2453 2407
rect 2462 2358 2466 2362
rect 2430 2338 2434 2342
rect 2478 2518 2482 2522
rect 2502 2548 2506 2552
rect 2478 2358 2482 2362
rect 2470 2308 2474 2312
rect 2442 2203 2446 2207
rect 2449 2203 2450 2207
rect 2450 2203 2453 2207
rect 2438 2068 2442 2072
rect 2442 2003 2446 2007
rect 2449 2003 2450 2007
rect 2450 2003 2453 2007
rect 2478 1868 2482 1872
rect 2442 1803 2446 1807
rect 2449 1803 2450 1807
rect 2450 1803 2453 1807
rect 2462 1758 2466 1762
rect 2442 1603 2446 1607
rect 2449 1603 2450 1607
rect 2450 1603 2453 1607
rect 2422 1508 2426 1512
rect 2398 1468 2402 1472
rect 2414 1468 2418 1472
rect 2442 1403 2446 1407
rect 2449 1403 2450 1407
rect 2450 1403 2453 1407
rect 2414 1288 2418 1292
rect 2358 1078 2362 1082
rect 2430 1308 2434 1312
rect 2442 1203 2446 1207
rect 2449 1203 2450 1207
rect 2450 1203 2453 1207
rect 2366 1048 2370 1052
rect 2406 1028 2410 1032
rect 2390 898 2394 902
rect 2318 868 2322 872
rect 2206 668 2210 672
rect 2358 718 2362 722
rect 2318 668 2322 672
rect 2174 578 2178 582
rect 2206 558 2210 562
rect 2078 148 2082 152
rect 2118 218 2122 222
rect 2126 158 2130 162
rect 2094 128 2098 132
rect 2054 68 2058 72
rect 1422 18 1426 22
rect 2086 18 2090 22
rect 2262 508 2266 512
rect 2318 448 2322 452
rect 2214 178 2218 182
rect 2222 148 2226 152
rect 2334 378 2338 382
rect 2270 288 2274 292
rect 2262 198 2266 202
rect 2286 188 2290 192
rect 2326 188 2330 192
rect 2442 1003 2446 1007
rect 2449 1003 2450 1007
rect 2450 1003 2453 1007
rect 2398 768 2402 772
rect 2442 803 2446 807
rect 2449 803 2450 807
rect 2450 803 2453 807
rect 2406 708 2410 712
rect 2390 438 2394 442
rect 2398 398 2402 402
rect 2414 648 2418 652
rect 2422 648 2426 652
rect 2442 603 2446 607
rect 2449 603 2450 607
rect 2450 603 2453 607
rect 2422 598 2426 602
rect 2502 2268 2506 2272
rect 2534 2528 2538 2532
rect 2534 2238 2538 2242
rect 2574 2358 2578 2362
rect 2590 2718 2594 2722
rect 2598 2478 2602 2482
rect 2582 2348 2586 2352
rect 2558 2148 2562 2152
rect 2526 2058 2530 2062
rect 2550 1988 2554 1992
rect 2510 1778 2514 1782
rect 2478 1378 2482 1382
rect 2510 1248 2514 1252
rect 2526 1388 2530 1392
rect 2582 2128 2586 2132
rect 3022 3028 3026 3032
rect 2806 2948 2810 2952
rect 2870 2948 2874 2952
rect 2910 2928 2914 2932
rect 2750 2908 2754 2912
rect 2750 2878 2754 2882
rect 2878 2888 2882 2892
rect 2654 2738 2658 2742
rect 2622 2718 2626 2722
rect 2638 2528 2642 2532
rect 2638 2378 2642 2382
rect 2670 2658 2674 2662
rect 2742 2748 2746 2752
rect 2686 2528 2690 2532
rect 2678 2478 2682 2482
rect 2678 2358 2682 2362
rect 2670 2348 2674 2352
rect 2694 2318 2698 2322
rect 2702 2308 2706 2312
rect 2638 2038 2642 2042
rect 2630 2018 2634 2022
rect 2606 1958 2610 1962
rect 2630 1958 2634 1962
rect 2590 1658 2594 1662
rect 2598 1548 2602 1552
rect 2566 1538 2570 1542
rect 2574 1538 2578 1542
rect 2678 2088 2682 2092
rect 2718 2088 2722 2092
rect 2694 2068 2698 2072
rect 2766 2658 2770 2662
rect 2774 2458 2778 2462
rect 2814 2748 2818 2752
rect 2910 2748 2914 2752
rect 2918 2648 2922 2652
rect 2798 2368 2802 2372
rect 2758 2278 2762 2282
rect 2750 2068 2754 2072
rect 2734 1998 2738 2002
rect 2742 1988 2746 1992
rect 2766 1918 2770 1922
rect 2822 2608 2826 2612
rect 2830 2388 2834 2392
rect 2798 2128 2802 2132
rect 2782 2058 2786 2062
rect 2798 1998 2802 2002
rect 2782 1958 2786 1962
rect 2790 1778 2794 1782
rect 2654 1698 2658 1702
rect 2622 1538 2626 1542
rect 2526 1288 2530 1292
rect 2534 1268 2538 1272
rect 2566 1158 2570 1162
rect 2518 1048 2522 1052
rect 2510 958 2514 962
rect 2502 938 2506 942
rect 2486 738 2490 742
rect 2462 428 2466 432
rect 2414 348 2418 352
rect 2382 268 2386 272
rect 2442 403 2446 407
rect 2449 403 2450 407
rect 2450 403 2453 407
rect 2494 388 2498 392
rect 2422 298 2426 302
rect 2414 258 2418 262
rect 2442 203 2446 207
rect 2449 203 2450 207
rect 2450 203 2453 207
rect 2422 138 2426 142
rect 2494 128 2498 132
rect 2174 28 2178 32
rect 2526 878 2530 882
rect 2510 728 2514 732
rect 2518 728 2522 732
rect 2526 718 2530 722
rect 2550 1058 2554 1062
rect 2558 978 2562 982
rect 2582 878 2586 882
rect 2638 1308 2642 1312
rect 2638 1128 2642 1132
rect 2630 958 2634 962
rect 2622 848 2626 852
rect 2542 808 2546 812
rect 2566 808 2570 812
rect 2534 508 2538 512
rect 2518 448 2522 452
rect 2534 448 2538 452
rect 2518 398 2522 402
rect 2534 378 2538 382
rect 2598 728 2602 732
rect 2590 658 2594 662
rect 2622 658 2626 662
rect 2614 558 2618 562
rect 2566 328 2570 332
rect 2534 178 2538 182
rect 2566 128 2570 132
rect 2606 68 2610 72
rect 2734 1688 2738 1692
rect 2750 1688 2754 1692
rect 2726 1468 2730 1472
rect 2734 1268 2738 1272
rect 2710 1238 2714 1242
rect 2654 1128 2658 1132
rect 2702 1118 2706 1122
rect 2734 1118 2738 1122
rect 2790 1588 2794 1592
rect 2782 1528 2786 1532
rect 2774 1268 2778 1272
rect 2838 2218 2842 2222
rect 2830 2148 2834 2152
rect 2830 2138 2834 2142
rect 2830 2088 2834 2092
rect 2814 1878 2818 1882
rect 2954 2903 2958 2907
rect 2961 2903 2962 2907
rect 2962 2903 2965 2907
rect 2954 2703 2958 2707
rect 2961 2703 2962 2707
rect 2962 2703 2965 2707
rect 2998 2738 3002 2742
rect 2990 2718 2994 2722
rect 3006 2558 3010 2562
rect 2954 2503 2958 2507
rect 2961 2503 2962 2507
rect 2962 2503 2965 2507
rect 2998 2478 3002 2482
rect 2954 2303 2958 2307
rect 2961 2303 2962 2307
rect 2962 2303 2965 2307
rect 3014 2298 3018 2302
rect 2990 2168 2994 2172
rect 2954 2103 2958 2107
rect 2961 2103 2962 2107
rect 2962 2103 2965 2107
rect 2942 1948 2946 1952
rect 2954 1903 2958 1907
rect 2961 1903 2962 1907
rect 2962 1903 2965 1907
rect 2974 1898 2978 1902
rect 3006 1838 3010 1842
rect 2954 1703 2958 1707
rect 2961 1703 2962 1707
rect 2962 1703 2965 1707
rect 2870 1638 2874 1642
rect 2878 1638 2882 1642
rect 2830 1628 2834 1632
rect 2822 1538 2826 1542
rect 2830 1518 2834 1522
rect 2798 1318 2802 1322
rect 2790 1148 2794 1152
rect 2670 878 2674 882
rect 2670 828 2674 832
rect 2662 768 2666 772
rect 2654 758 2658 762
rect 2678 738 2682 742
rect 2694 728 2698 732
rect 2678 588 2682 592
rect 2662 128 2666 132
rect 2678 478 2682 482
rect 2774 1058 2778 1062
rect 2750 1008 2754 1012
rect 2710 808 2714 812
rect 2726 758 2730 762
rect 2718 718 2722 722
rect 2726 658 2730 662
rect 2702 148 2706 152
rect 2694 128 2698 132
rect 2718 78 2722 82
rect 2774 868 2778 872
rect 2766 838 2770 842
rect 2774 768 2778 772
rect 2822 1468 2826 1472
rect 2822 1128 2826 1132
rect 2774 558 2778 562
rect 2774 448 2778 452
rect 2854 1518 2858 1522
rect 2870 1488 2874 1492
rect 2846 1428 2850 1432
rect 2846 1328 2850 1332
rect 2838 1208 2842 1212
rect 2830 548 2834 552
rect 2870 1298 2874 1302
rect 2894 1458 2898 1462
rect 2886 1438 2890 1442
rect 2902 1218 2906 1222
rect 2886 1088 2890 1092
rect 2878 1008 2882 1012
rect 2886 898 2890 902
rect 2886 878 2890 882
rect 2894 828 2898 832
rect 2878 718 2882 722
rect 2886 708 2890 712
rect 2982 1578 2986 1582
rect 2942 1508 2946 1512
rect 2982 1508 2986 1512
rect 2954 1503 2958 1507
rect 2961 1503 2962 1507
rect 2962 1503 2965 1507
rect 2926 1298 2930 1302
rect 2954 1303 2958 1307
rect 2961 1303 2962 1307
rect 2962 1303 2965 1307
rect 2974 1298 2978 1302
rect 2954 1103 2958 1107
rect 2961 1103 2962 1107
rect 2962 1103 2965 1107
rect 3014 1458 3018 1462
rect 3014 1128 3018 1132
rect 3006 1118 3010 1122
rect 2998 1108 3002 1112
rect 2982 1088 2986 1092
rect 3014 1088 3018 1092
rect 2942 1048 2946 1052
rect 2998 1038 3002 1042
rect 2998 1008 3002 1012
rect 3342 2958 3346 2962
rect 3062 2658 3066 2662
rect 3030 2288 3034 2292
rect 3038 2288 3042 2292
rect 3062 2078 3066 2082
rect 3358 2868 3362 2872
rect 3190 2728 3194 2732
rect 3190 2658 3194 2662
rect 3078 2348 3082 2352
rect 3086 2278 3090 2282
rect 3126 2238 3130 2242
rect 3102 2078 3106 2082
rect 3150 2268 3154 2272
rect 3238 2548 3242 2552
rect 3222 2538 3226 2542
rect 3270 2528 3274 2532
rect 3254 2518 3258 2522
rect 3206 2468 3210 2472
rect 3166 2338 3170 2342
rect 3078 1958 3082 1962
rect 3078 1938 3082 1942
rect 3142 1938 3146 1942
rect 3150 1938 3154 1942
rect 3206 2348 3210 2352
rect 3238 2338 3242 2342
rect 3086 1708 3090 1712
rect 3110 1718 3114 1722
rect 3094 1618 3098 1622
rect 3102 1618 3106 1622
rect 3102 1558 3106 1562
rect 3134 1728 3138 1732
rect 3158 1648 3162 1652
rect 3166 1648 3170 1652
rect 3182 1628 3186 1632
rect 3118 1508 3122 1512
rect 3110 1448 3114 1452
rect 3070 1228 3074 1232
rect 3062 1188 3066 1192
rect 3062 1158 3066 1162
rect 3062 1018 3066 1022
rect 2954 903 2958 907
rect 2961 903 2962 907
rect 2962 903 2965 907
rect 2942 868 2946 872
rect 2934 858 2938 862
rect 2918 818 2922 822
rect 2894 628 2898 632
rect 2974 818 2978 822
rect 2954 703 2958 707
rect 2961 703 2962 707
rect 2962 703 2965 707
rect 2926 648 2930 652
rect 2918 618 2922 622
rect 2954 503 2958 507
rect 2961 503 2962 507
rect 2962 503 2965 507
rect 2950 488 2954 492
rect 3006 648 3010 652
rect 2926 438 2930 442
rect 2894 348 2898 352
rect 2806 278 2810 282
rect 2926 328 2930 332
rect 2934 298 2938 302
rect 2854 248 2858 252
rect 2954 303 2958 307
rect 2961 303 2962 307
rect 2962 303 2965 307
rect 2998 508 3002 512
rect 3006 448 3010 452
rect 3102 1158 3106 1162
rect 3110 1138 3114 1142
rect 3086 1078 3090 1082
rect 3110 1078 3114 1082
rect 3086 1038 3090 1042
rect 3070 938 3074 942
rect 3126 978 3130 982
rect 3166 1578 3170 1582
rect 3238 2178 3242 2182
rect 3230 2148 3234 2152
rect 3214 2138 3218 2142
rect 3270 2188 3274 2192
rect 3254 2078 3258 2082
rect 3222 1998 3226 2002
rect 3214 1948 3218 1952
rect 3254 1938 3258 1942
rect 3326 2458 3330 2462
rect 3302 2268 3306 2272
rect 3302 2048 3306 2052
rect 3366 2418 3370 2422
rect 3350 2278 3354 2282
rect 3342 2258 3346 2262
rect 3474 3003 3478 3007
rect 3481 3003 3482 3007
rect 3482 3003 3485 3007
rect 3398 2928 3402 2932
rect 3390 2918 3394 2922
rect 3474 2803 3478 2807
rect 3481 2803 3482 2807
rect 3482 2803 3485 2807
rect 3470 2768 3474 2772
rect 3430 2748 3434 2752
rect 3390 2548 3394 2552
rect 3710 2938 3714 2942
rect 3510 2738 3514 2742
rect 3474 2603 3478 2607
rect 3481 2603 3482 2607
rect 3482 2603 3485 2607
rect 3590 2868 3594 2872
rect 3590 2688 3594 2692
rect 3422 2528 3426 2532
rect 3398 2278 3402 2282
rect 3374 2258 3378 2262
rect 3334 2048 3338 2052
rect 3350 1948 3354 1952
rect 3214 1758 3218 1762
rect 3246 1648 3250 1652
rect 3214 1628 3218 1632
rect 3206 1548 3210 1552
rect 3150 1528 3154 1532
rect 3174 1528 3178 1532
rect 3238 1538 3242 1542
rect 3222 1478 3226 1482
rect 3198 1218 3202 1222
rect 3206 1158 3210 1162
rect 3150 1118 3154 1122
rect 3150 988 3154 992
rect 3134 958 3138 962
rect 3118 898 3122 902
rect 3086 888 3090 892
rect 3102 888 3106 892
rect 3198 1018 3202 1022
rect 3078 808 3082 812
rect 3134 788 3138 792
rect 3110 738 3114 742
rect 2954 103 2958 107
rect 2961 103 2962 107
rect 2962 103 2965 107
rect 2974 88 2978 92
rect 3094 478 3098 482
rect 3118 478 3122 482
rect 3094 448 3098 452
rect 3118 438 3122 442
rect 3158 708 3162 712
rect 3190 858 3194 862
rect 3182 838 3186 842
rect 3198 828 3202 832
rect 3198 638 3202 642
rect 3302 1648 3306 1652
rect 3310 1588 3314 1592
rect 3318 1558 3322 1562
rect 3366 1548 3370 1552
rect 3310 1478 3314 1482
rect 3294 1468 3298 1472
rect 3350 1538 3354 1542
rect 3334 1528 3338 1532
rect 3374 1528 3378 1532
rect 3526 2458 3530 2462
rect 3542 2458 3546 2462
rect 3502 2438 3506 2442
rect 3474 2403 3478 2407
rect 3481 2403 3482 2407
rect 3482 2403 3485 2407
rect 3422 2248 3426 2252
rect 3414 2068 3418 2072
rect 3406 2058 3410 2062
rect 3474 2203 3478 2207
rect 3481 2203 3482 2207
rect 3482 2203 3485 2207
rect 3574 2238 3578 2242
rect 3518 2068 3522 2072
rect 3474 2003 3478 2007
rect 3481 2003 3482 2007
rect 3482 2003 3485 2007
rect 3414 1748 3418 1752
rect 3390 1698 3394 1702
rect 3382 1458 3386 1462
rect 3326 1448 3330 1452
rect 3374 1448 3378 1452
rect 3254 1268 3258 1272
rect 3254 1258 3258 1262
rect 3246 1238 3250 1242
rect 3238 1218 3242 1222
rect 3230 1128 3234 1132
rect 3254 1138 3258 1142
rect 3286 1318 3290 1322
rect 3342 1338 3346 1342
rect 3358 1338 3362 1342
rect 3310 1308 3314 1312
rect 3262 1058 3266 1062
rect 3326 1308 3330 1312
rect 3302 928 3306 932
rect 3310 918 3314 922
rect 3318 898 3322 902
rect 3230 678 3234 682
rect 3262 698 3266 702
rect 3246 668 3250 672
rect 3238 588 3242 592
rect 3214 558 3218 562
rect 3182 488 3186 492
rect 3142 288 3146 292
rect 3246 528 3250 532
rect 3230 508 3234 512
rect 3262 398 3266 402
rect 3230 378 3234 382
rect 3254 358 3258 362
rect 3302 788 3306 792
rect 3302 688 3306 692
rect 3366 1238 3370 1242
rect 3334 1048 3338 1052
rect 3350 918 3354 922
rect 3366 768 3370 772
rect 3398 1558 3402 1562
rect 3422 1468 3426 1472
rect 3474 1803 3478 1807
rect 3481 1803 3482 1807
rect 3482 1803 3485 1807
rect 3526 1898 3530 1902
rect 3518 1848 3522 1852
rect 3526 1768 3530 1772
rect 3446 1678 3450 1682
rect 3422 1298 3426 1302
rect 3438 1268 3442 1272
rect 3446 1188 3450 1192
rect 3486 1678 3490 1682
rect 3470 1638 3474 1642
rect 3474 1603 3478 1607
rect 3481 1603 3482 1607
rect 3482 1603 3485 1607
rect 3502 1538 3506 1542
rect 3670 2878 3674 2882
rect 3630 2728 3634 2732
rect 3654 2688 3658 2692
rect 3606 2588 3610 2592
rect 3622 2488 3626 2492
rect 3694 2568 3698 2572
rect 3654 2428 3658 2432
rect 3654 2238 3658 2242
rect 3582 1558 3586 1562
rect 3542 1548 3546 1552
rect 3526 1528 3530 1532
rect 3470 1508 3474 1512
rect 3474 1403 3478 1407
rect 3481 1403 3482 1407
rect 3482 1403 3485 1407
rect 3474 1203 3478 1207
rect 3481 1203 3482 1207
rect 3482 1203 3485 1207
rect 3486 1148 3490 1152
rect 3542 1488 3546 1492
rect 3502 1308 3506 1312
rect 3542 1348 3546 1352
rect 3646 1978 3650 1982
rect 3630 1758 3634 1762
rect 3654 1758 3658 1762
rect 3622 1418 3626 1422
rect 3558 1168 3562 1172
rect 3446 1078 3450 1082
rect 3470 1048 3474 1052
rect 3526 1038 3530 1042
rect 3474 1003 3478 1007
rect 3481 1003 3482 1007
rect 3482 1003 3485 1007
rect 3414 928 3418 932
rect 3422 918 3426 922
rect 3398 858 3402 862
rect 3366 658 3370 662
rect 3294 528 3298 532
rect 3310 458 3314 462
rect 3326 408 3330 412
rect 3422 708 3426 712
rect 3430 698 3434 702
rect 3390 688 3394 692
rect 3502 818 3506 822
rect 3474 803 3478 807
rect 3481 803 3482 807
rect 3482 803 3485 807
rect 3406 298 3410 302
rect 3510 718 3514 722
rect 3502 678 3506 682
rect 3474 603 3478 607
rect 3481 603 3482 607
rect 3482 603 3485 607
rect 3474 403 3478 407
rect 3481 403 3482 407
rect 3482 403 3485 407
rect 3454 238 3458 242
rect 3470 238 3474 242
rect 3422 228 3426 232
rect 3590 1058 3594 1062
rect 3590 928 3594 932
rect 3542 668 3546 672
rect 3566 788 3570 792
rect 3622 1318 3626 1322
rect 3622 1258 3626 1262
rect 3622 1188 3626 1192
rect 3622 938 3626 942
rect 3646 1348 3650 1352
rect 3758 2738 3762 2742
rect 3742 2638 3746 2642
rect 3798 2768 3802 2772
rect 3710 2128 3714 2132
rect 3742 2228 3746 2232
rect 3838 2718 3842 2722
rect 3830 2528 3834 2532
rect 3814 2338 3818 2342
rect 3902 2358 3906 2362
rect 3870 2328 3874 2332
rect 3854 2298 3858 2302
rect 3782 2148 3786 2152
rect 3822 2078 3826 2082
rect 3862 2188 3866 2192
rect 3918 2288 3922 2292
rect 3978 2903 3982 2907
rect 3985 2903 3986 2907
rect 3986 2903 3989 2907
rect 3958 2748 3962 2752
rect 4062 2748 4066 2752
rect 4102 2748 4106 2752
rect 3998 2728 4002 2732
rect 4094 2728 4098 2732
rect 3978 2703 3982 2707
rect 3985 2703 3986 2707
rect 3986 2703 3989 2707
rect 4086 2688 4090 2692
rect 4038 2628 4042 2632
rect 3978 2503 3982 2507
rect 3985 2503 3986 2507
rect 3986 2503 3989 2507
rect 3978 2303 3982 2307
rect 3985 2303 3986 2307
rect 3986 2303 3989 2307
rect 4126 2958 4130 2962
rect 4150 2958 4154 2962
rect 4126 2738 4130 2742
rect 4054 2488 4058 2492
rect 3982 2278 3986 2282
rect 3894 2068 3898 2072
rect 3806 2058 3810 2062
rect 3766 1968 3770 1972
rect 3710 1858 3714 1862
rect 3702 1788 3706 1792
rect 3694 1668 3698 1672
rect 3694 1528 3698 1532
rect 3670 1338 3674 1342
rect 3694 1278 3698 1282
rect 3750 1888 3754 1892
rect 3758 1858 3762 1862
rect 3758 1738 3762 1742
rect 3750 1668 3754 1672
rect 3766 1528 3770 1532
rect 3726 1218 3730 1222
rect 3710 1178 3714 1182
rect 3686 858 3690 862
rect 3638 728 3642 732
rect 3526 318 3530 322
rect 3710 1058 3714 1062
rect 3790 1708 3794 1712
rect 3774 1268 3778 1272
rect 3758 1258 3762 1262
rect 3822 1848 3826 1852
rect 3830 1698 3834 1702
rect 3830 1558 3834 1562
rect 3830 1548 3834 1552
rect 3782 1168 3786 1172
rect 3758 1128 3762 1132
rect 3734 1068 3738 1072
rect 3758 938 3762 942
rect 3766 928 3770 932
rect 3710 688 3714 692
rect 3702 658 3706 662
rect 3870 1288 3874 1292
rect 3918 1758 3922 1762
rect 3926 1618 3930 1622
rect 3934 1578 3938 1582
rect 3950 1678 3954 1682
rect 3950 1568 3954 1572
rect 3878 1278 3882 1282
rect 3830 1048 3834 1052
rect 3814 1028 3818 1032
rect 3814 938 3818 942
rect 3806 738 3810 742
rect 3726 508 3730 512
rect 3670 438 3674 442
rect 3702 358 3706 362
rect 3686 298 3690 302
rect 3474 203 3478 207
rect 3481 203 3482 207
rect 3482 203 3485 207
rect 3574 178 3578 182
rect 3454 168 3458 172
rect 3182 128 3186 132
rect 3350 118 3354 122
rect 3174 68 3178 72
rect 3638 178 3642 182
rect 3726 338 3730 342
rect 3726 318 3730 322
rect 3750 348 3754 352
rect 3886 1128 3890 1132
rect 3958 1108 3962 1112
rect 3958 1058 3962 1062
rect 3902 838 3906 842
rect 3830 148 3834 152
rect 3854 368 3858 372
rect 3878 668 3882 672
rect 3958 888 3962 892
rect 3926 868 3930 872
rect 3934 748 3938 752
rect 3902 578 3906 582
rect 3934 538 3938 542
rect 3902 518 3906 522
rect 3894 448 3898 452
rect 3886 328 3890 332
rect 3886 308 3890 312
rect 3910 358 3914 362
rect 3902 238 3906 242
rect 3942 368 3946 372
rect 3978 2103 3982 2107
rect 3985 2103 3986 2107
rect 3986 2103 3989 2107
rect 3998 1948 4002 1952
rect 3978 1903 3982 1907
rect 3985 1903 3986 1907
rect 3986 1903 3989 1907
rect 3978 1703 3982 1707
rect 3985 1703 3986 1707
rect 3986 1703 3989 1707
rect 3978 1503 3982 1507
rect 3985 1503 3986 1507
rect 3986 1503 3989 1507
rect 4022 2068 4026 2072
rect 4030 2038 4034 2042
rect 4046 2078 4050 2082
rect 4006 1848 4010 1852
rect 4038 1818 4042 1822
rect 4078 2158 4082 2162
rect 4078 2098 4082 2102
rect 4062 2078 4066 2082
rect 4070 2068 4074 2072
rect 4054 1748 4058 1752
rect 4030 1728 4034 1732
rect 4046 1518 4050 1522
rect 3998 1438 4002 1442
rect 4014 1378 4018 1382
rect 4046 1368 4050 1372
rect 3978 1303 3982 1307
rect 3985 1303 3986 1307
rect 3986 1303 3989 1307
rect 4014 1268 4018 1272
rect 3998 1148 4002 1152
rect 3978 1103 3982 1107
rect 3985 1103 3986 1107
rect 3986 1103 3989 1107
rect 3998 928 4002 932
rect 3978 903 3982 907
rect 3985 903 3986 907
rect 3986 903 3989 907
rect 4006 728 4010 732
rect 3978 703 3982 707
rect 3985 703 3986 707
rect 3986 703 3989 707
rect 3978 503 3982 507
rect 3985 503 3986 507
rect 3986 503 3989 507
rect 3998 468 4002 472
rect 3998 418 4002 422
rect 3958 328 3962 332
rect 3974 318 3978 322
rect 3978 303 3982 307
rect 3985 303 3986 307
rect 3986 303 3989 307
rect 3966 278 3970 282
rect 3978 103 3982 107
rect 3985 103 3986 107
rect 3986 103 3989 107
rect 3590 68 3594 72
rect 3686 68 3690 72
rect 4030 328 4034 332
rect 4054 1248 4058 1252
rect 4054 748 4058 752
rect 4150 2258 4154 2262
rect 4102 2138 4106 2142
rect 4118 2078 4122 2082
rect 4110 1868 4114 1872
rect 4094 1438 4098 1442
rect 4078 668 4082 672
rect 4078 568 4082 572
rect 4070 558 4074 562
rect 4078 388 4082 392
rect 4078 268 4082 272
rect 4070 258 4074 262
rect 4070 228 4074 232
rect 4062 218 4066 222
rect 4118 1648 4122 1652
rect 4142 1888 4146 1892
rect 4142 1688 4146 1692
rect 4126 1358 4130 1362
rect 4150 1328 4154 1332
rect 4166 2488 4170 2492
rect 4174 1928 4178 1932
rect 4166 1758 4170 1762
rect 4174 1538 4178 1542
rect 4190 2938 4194 2942
rect 4254 3068 4258 3072
rect 4230 3058 4234 3062
rect 4270 3048 4274 3052
rect 4278 3038 4282 3042
rect 4302 3028 4306 3032
rect 4214 2948 4218 2952
rect 4246 2768 4250 2772
rect 4238 2748 4242 2752
rect 4238 2738 4242 2742
rect 4222 2578 4226 2582
rect 4190 1568 4194 1572
rect 4110 878 4114 882
rect 4102 758 4106 762
rect 4110 528 4114 532
rect 4142 1058 4146 1062
rect 4166 1048 4170 1052
rect 4174 278 4178 282
rect 4174 108 4178 112
rect 4150 98 4154 102
rect 4142 78 4146 82
rect 3726 58 3730 62
rect 4262 2428 4266 2432
rect 4238 2028 4242 2032
rect 4230 1698 4234 1702
rect 4230 1468 4234 1472
rect 4254 1748 4258 1752
rect 4246 1708 4250 1712
rect 4222 1288 4226 1292
rect 4222 1088 4226 1092
rect 4222 1018 4226 1022
rect 4222 1008 4226 1012
rect 4214 968 4218 972
rect 4206 878 4210 882
rect 4206 778 4210 782
rect 4262 1468 4266 1472
rect 4246 1048 4250 1052
rect 4238 1038 4242 1042
rect 4246 948 4250 952
rect 4270 1018 4274 1022
rect 4254 778 4258 782
rect 4294 2748 4298 2752
rect 4294 2268 4298 2272
rect 4286 1798 4290 1802
rect 4350 3058 4354 3062
rect 4334 2748 4338 2752
rect 4326 2738 4330 2742
rect 4318 2348 4322 2352
rect 4302 1728 4306 1732
rect 4286 1238 4290 1242
rect 4286 1168 4290 1172
rect 4238 288 4242 292
rect 4286 348 4290 352
rect 4206 188 4210 192
rect 4310 848 4314 852
rect 4302 638 4306 642
rect 4294 158 4298 162
rect 4302 148 4306 152
rect 4302 138 4306 142
rect 4198 88 4202 92
rect 4342 2648 4346 2652
rect 4326 2098 4330 2102
rect 4366 2448 4370 2452
rect 4366 2428 4370 2432
rect 4334 1828 4338 1832
rect 4334 1798 4338 1802
rect 4342 1788 4346 1792
rect 4342 1778 4346 1782
rect 4334 1118 4338 1122
rect 4382 2368 4386 2372
rect 4350 1108 4354 1112
rect 4358 1088 4362 1092
rect 4342 478 4346 482
rect 4326 448 4330 452
rect 4366 158 4370 162
rect 4326 128 4330 132
rect 4318 68 4322 72
rect 4174 38 4178 42
rect 394 3 398 7
rect 401 3 402 7
rect 402 3 405 7
rect 1418 3 1422 7
rect 1425 3 1426 7
rect 1426 3 1429 7
rect 2442 3 2446 7
rect 2449 3 2450 7
rect 2450 3 2453 7
rect 3474 3 3478 7
rect 3481 3 3482 7
rect 3482 3 3485 7
<< metal5 >>
rect 902 3103 905 3107
rect 901 3102 906 3103
rect 911 3102 912 3107
rect 1934 3103 1937 3107
rect 1933 3102 1938 3103
rect 1943 3102 1944 3107
rect 2958 3103 2961 3107
rect 2957 3102 2962 3103
rect 2967 3102 2968 3107
rect 3982 3103 3985 3107
rect 3981 3102 3986 3103
rect 3991 3102 3992 3107
rect 226 3068 630 3071
rect 4258 3068 4301 3071
rect 322 3058 702 3061
rect 4234 3058 4350 3061
rect 4258 3048 4270 3051
rect 4274 3038 4278 3041
rect 3026 3028 4302 3031
rect 398 3003 401 3007
rect 397 3002 402 3003
rect 407 3002 408 3007
rect 1422 3003 1425 3007
rect 1421 3002 1426 3003
rect 1431 3002 1432 3007
rect 2446 3003 2449 3007
rect 2445 3002 2450 3003
rect 2455 3002 2456 3007
rect 3478 3003 3481 3007
rect 3477 3002 3482 3003
rect 3487 3002 3488 3007
rect 3346 2958 4126 2961
rect 1466 2948 1678 2951
rect 2810 2948 2870 2951
rect 4150 2951 4153 2958
rect 4150 2948 4214 2951
rect 3714 2938 4190 2941
rect 2914 2928 3398 2931
rect 2418 2918 3390 2921
rect 1986 2908 2750 2911
rect 902 2903 905 2907
rect 901 2902 906 2903
rect 911 2902 912 2907
rect 1934 2903 1937 2907
rect 1933 2902 1938 2903
rect 1943 2902 1944 2907
rect 2958 2903 2961 2907
rect 2957 2902 2962 2903
rect 2967 2902 2968 2907
rect 3982 2903 3985 2907
rect 3981 2902 3986 2903
rect 3991 2902 3992 2907
rect 1602 2888 2878 2891
rect 1754 2878 2158 2881
rect 2754 2878 3670 2881
rect 1562 2868 2446 2871
rect 3362 2868 3590 2871
rect 398 2803 401 2807
rect 397 2802 402 2803
rect 407 2802 408 2807
rect 1422 2803 1425 2807
rect 1421 2802 1426 2803
rect 1431 2802 1432 2807
rect 2446 2803 2449 2807
rect 2445 2802 2450 2803
rect 2455 2802 2456 2807
rect 3478 2803 3481 2807
rect 3477 2802 3482 2803
rect 3487 2802 3488 2807
rect 3474 2768 3798 2771
rect 4130 2768 4246 2771
rect 3202 2758 4297 2761
rect 4294 2752 4297 2758
rect 802 2748 1006 2751
rect 2746 2748 2814 2751
rect 2914 2748 3430 2751
rect 3962 2748 4062 2751
rect 4106 2748 4238 2751
rect 4338 2748 4349 2751
rect 2226 2738 2654 2741
rect 2658 2738 2998 2741
rect 3514 2738 3758 2741
rect 4118 2738 4126 2741
rect 4130 2738 4238 2741
rect 4322 2738 4326 2741
rect 2322 2728 3190 2731
rect 3634 2728 3998 2731
rect 2594 2718 2622 2721
rect 2626 2718 2990 2721
rect 4094 2721 4097 2728
rect 3842 2718 4097 2721
rect 902 2703 905 2707
rect 901 2702 906 2703
rect 911 2702 912 2707
rect 1934 2703 1937 2707
rect 1933 2702 1938 2703
rect 1943 2702 1944 2707
rect 2958 2703 2961 2707
rect 2957 2702 2962 2703
rect 2967 2702 2968 2707
rect 3982 2703 3985 2707
rect 3981 2702 3986 2703
rect 3991 2702 3992 2707
rect 2098 2688 3590 2691
rect 3658 2688 4086 2691
rect 1986 2658 2670 2661
rect 2674 2658 2766 2661
rect 3066 2658 3190 2661
rect 2098 2648 2918 2651
rect 4306 2648 4342 2651
rect 1898 2638 3742 2641
rect 1290 2628 4038 2631
rect 2050 2618 2825 2621
rect 2822 2612 2825 2618
rect 398 2603 401 2607
rect 397 2602 402 2603
rect 407 2602 408 2607
rect 1422 2603 1425 2607
rect 1421 2602 1426 2603
rect 1431 2602 1432 2607
rect 2446 2603 2449 2607
rect 2445 2602 2450 2603
rect 2455 2602 2456 2607
rect 3478 2603 3481 2607
rect 3477 2602 3482 2603
rect 3487 2602 3488 2607
rect 1754 2588 3606 2591
rect 2090 2578 4222 2581
rect 2018 2568 3694 2571
rect 122 2558 574 2561
rect 2266 2558 3006 2561
rect 1818 2548 2502 2551
rect 3242 2548 3390 2551
rect 2426 2538 3222 2541
rect 1510 2531 1513 2538
rect 834 2528 1806 2531
rect 1866 2528 2086 2531
rect 2538 2528 2638 2531
rect 2690 2528 3270 2531
rect 3426 2528 3830 2531
rect 2482 2518 3254 2521
rect 902 2503 905 2507
rect 901 2502 906 2503
rect 911 2502 912 2507
rect 1934 2503 1937 2507
rect 1933 2502 1938 2503
rect 1943 2502 1944 2507
rect 2958 2503 2961 2507
rect 2957 2502 2962 2503
rect 2967 2502 2968 2507
rect 3982 2503 3985 2507
rect 3981 2502 3986 2503
rect 3991 2502 3992 2507
rect 1954 2498 2294 2501
rect 2362 2498 2941 2501
rect 1810 2488 3622 2491
rect 4058 2488 4166 2491
rect 1682 2478 1734 2481
rect 1922 2478 2598 2481
rect 2682 2478 2998 2481
rect 2946 2468 3101 2471
rect 3106 2468 3206 2471
rect 826 2458 1374 2461
rect 1378 2458 1678 2461
rect 1858 2458 2086 2461
rect 2266 2458 2774 2461
rect 3330 2458 3526 2461
rect 3530 2458 3542 2461
rect 1362 2448 1446 2451
rect 1914 2448 2374 2451
rect 4366 2442 4369 2448
rect 1706 2438 2054 2441
rect 2178 2438 3502 2441
rect 1658 2428 1846 2431
rect 2002 2428 3654 2431
rect 4266 2428 4366 2431
rect 2226 2418 3366 2421
rect 1522 2408 2142 2411
rect 2146 2408 2358 2411
rect 398 2403 401 2407
rect 397 2402 402 2403
rect 407 2402 408 2407
rect 1422 2403 1425 2407
rect 1421 2402 1426 2403
rect 1431 2402 1432 2407
rect 2446 2403 2449 2407
rect 2445 2402 2450 2403
rect 2455 2402 2456 2407
rect 3478 2403 3481 2407
rect 3477 2402 3482 2403
rect 3487 2402 3488 2407
rect 1650 2388 2830 2391
rect 2426 2378 2638 2381
rect 1834 2368 2078 2371
rect 2410 2368 2798 2371
rect 4382 2362 4385 2368
rect 1762 2358 1982 2361
rect 2066 2358 2462 2361
rect 2482 2358 2574 2361
rect 2682 2358 3902 2361
rect 1402 2348 1766 2351
rect 1786 2348 1869 2351
rect 2098 2348 2182 2351
rect 2330 2348 2582 2351
rect 2586 2348 2670 2351
rect 3082 2348 3206 2351
rect 4306 2348 4318 2351
rect 1998 2342 2001 2347
rect 1122 2338 1846 2341
rect 2434 2338 3166 2341
rect 3242 2338 3814 2341
rect 2314 2328 3870 2331
rect 1090 2318 1622 2321
rect 1866 2318 1869 2321
rect 2234 2318 2694 2321
rect 2186 2308 2470 2311
rect 2474 2308 2702 2311
rect 902 2303 905 2307
rect 901 2302 906 2303
rect 911 2302 912 2307
rect 1934 2303 1937 2307
rect 1933 2302 1938 2303
rect 1943 2302 1944 2307
rect 2958 2303 2961 2307
rect 2957 2302 2962 2303
rect 2967 2302 2968 2307
rect 3982 2303 3985 2307
rect 3981 2302 3986 2303
rect 3991 2302 3992 2307
rect 2018 2298 2110 2301
rect 3018 2298 3854 2301
rect 1858 2288 1966 2291
rect 2226 2288 3030 2291
rect 3042 2288 3918 2291
rect 1706 2278 2014 2281
rect 2762 2278 3086 2281
rect 3090 2278 3350 2281
rect 3402 2278 3982 2281
rect 1338 2268 1606 2271
rect 2394 2268 2502 2271
rect 3154 2268 3302 2271
rect 818 2258 838 2261
rect 1042 2258 1718 2261
rect 1850 2258 2126 2261
rect 3346 2258 3374 2261
rect 4294 2261 4297 2268
rect 4154 2258 4297 2261
rect 1866 2248 1990 2251
rect 2010 2248 2022 2251
rect 2298 2248 3422 2251
rect 1990 2241 1993 2248
rect 1990 2238 2534 2241
rect 3130 2238 3574 2241
rect 3578 2238 3654 2241
rect 1802 2228 1982 2231
rect 2410 2228 3742 2231
rect 2290 2218 2838 2221
rect 398 2203 401 2207
rect 397 2202 402 2203
rect 407 2202 408 2207
rect 1422 2203 1425 2207
rect 1421 2202 1426 2203
rect 1431 2202 1432 2207
rect 2446 2203 2449 2207
rect 2445 2202 2450 2203
rect 2455 2202 2456 2207
rect 3478 2203 3481 2207
rect 3477 2202 3482 2203
rect 3487 2202 3488 2207
rect 1998 2188 3270 2191
rect 1998 2181 2001 2188
rect 3282 2188 3862 2191
rect 1762 2178 2001 2181
rect 2010 2178 3238 2181
rect 186 2168 1766 2171
rect 2058 2168 2990 2171
rect 810 2158 838 2161
rect 1530 2158 2254 2161
rect 4078 2152 4081 2158
rect 34 2148 190 2151
rect 850 2148 918 2151
rect 1810 2148 2294 2151
rect 2562 2148 2830 2151
rect 3234 2148 3782 2151
rect 4098 2148 4105 2151
rect 4102 2142 4105 2148
rect 818 2138 902 2141
rect 906 2138 1014 2141
rect 2002 2138 2257 2141
rect 2834 2138 3214 2141
rect 2254 2132 2257 2138
rect 2306 2128 2582 2131
rect 2802 2128 3710 2131
rect 902 2103 905 2107
rect 901 2102 906 2103
rect 911 2102 912 2107
rect 1934 2103 1937 2107
rect 1933 2102 1938 2103
rect 1943 2102 1944 2107
rect 2958 2103 2961 2107
rect 2957 2102 2962 2103
rect 2967 2102 2968 2107
rect 3982 2103 3985 2107
rect 3981 2102 3986 2103
rect 3991 2102 3992 2107
rect 1354 2098 1697 2101
rect 4082 2098 4326 2101
rect 1694 2092 1697 2098
rect 1842 2088 2214 2091
rect 2218 2088 2678 2091
rect 2722 2088 2830 2091
rect 646 2081 649 2088
rect 646 2078 1326 2081
rect 2346 2078 3062 2081
rect 3106 2078 3254 2081
rect 3826 2078 4046 2081
rect 4066 2078 4118 2081
rect 2442 2068 2694 2071
rect 2754 2068 3414 2071
rect 3522 2068 3894 2071
rect 4026 2068 4070 2071
rect 1726 2062 1729 2067
rect 650 2058 1070 2061
rect 2530 2058 2782 2061
rect 3410 2058 3806 2061
rect 530 2048 702 2051
rect 778 2048 1174 2051
rect 1642 2048 3277 2051
rect 3306 2048 3334 2051
rect 370 2038 1582 2041
rect 1874 2038 1950 2041
rect 2642 2038 4030 2041
rect 1322 2028 2062 2031
rect 4238 2022 4241 2028
rect 1970 2018 2630 2021
rect 1886 2011 1889 2018
rect 1834 2008 1889 2011
rect 398 2003 401 2007
rect 397 2002 402 2003
rect 407 2002 408 2007
rect 1422 2003 1425 2007
rect 1421 2002 1426 2003
rect 1431 2002 1432 2007
rect 2446 2003 2449 2007
rect 2445 2002 2450 2003
rect 2455 2002 2456 2007
rect 3478 2003 3481 2007
rect 3477 2002 3482 2003
rect 3487 2002 3488 2007
rect 2738 1998 2798 2001
rect 2802 1998 3222 2001
rect 1954 1988 2550 1991
rect 2554 1988 2742 1991
rect 1026 1978 1142 1981
rect 1466 1978 2142 1981
rect 2162 1978 3646 1981
rect 730 1968 998 1971
rect 1178 1968 1366 1971
rect 1370 1968 1750 1971
rect 1938 1968 3766 1971
rect 1138 1958 1750 1961
rect 2146 1958 2606 1961
rect 2610 1958 2630 1961
rect 2786 1958 3078 1961
rect 1586 1948 2166 1951
rect 2946 1948 3214 1951
rect 3354 1948 3998 1951
rect 162 1938 182 1941
rect 722 1938 918 1941
rect 1242 1938 1278 1941
rect 1906 1938 1910 1941
rect 3082 1938 3142 1941
rect 3154 1938 3254 1941
rect 4174 1938 4189 1941
rect 4174 1932 4177 1938
rect 194 1928 1142 1931
rect 1418 1928 1934 1931
rect 434 1918 1446 1921
rect 1506 1918 2766 1921
rect 1330 1908 1806 1911
rect 870 1901 873 1908
rect 902 1903 905 1907
rect 901 1902 906 1903
rect 911 1902 912 1907
rect 1934 1903 1937 1907
rect 1933 1902 1938 1903
rect 1943 1902 1944 1907
rect 2958 1903 2961 1907
rect 2957 1902 2962 1903
rect 2967 1902 2968 1907
rect 3982 1903 3985 1907
rect 3981 1902 3986 1903
rect 3991 1902 3992 1907
rect 682 1898 873 1901
rect 1138 1898 1574 1901
rect 2978 1898 3526 1901
rect 298 1888 822 1891
rect 842 1888 1118 1891
rect 1466 1888 1766 1891
rect 2058 1888 3750 1891
rect 538 1878 846 1881
rect 874 1878 1281 1881
rect 1290 1878 1718 1881
rect 4142 1881 4145 1888
rect 2818 1878 4145 1881
rect 394 1868 1134 1871
rect 1278 1871 1281 1878
rect 1278 1868 1510 1871
rect 1666 1868 1670 1871
rect 1674 1868 1718 1871
rect 2482 1868 4110 1871
rect 730 1858 998 1861
rect 1618 1858 1742 1861
rect 1762 1858 1894 1861
rect 1898 1858 2062 1861
rect 3714 1858 3758 1861
rect 2102 1851 2105 1858
rect 1378 1848 2105 1851
rect 3522 1848 3822 1851
rect 4002 1848 4006 1851
rect 1842 1838 3006 1841
rect 914 1828 1454 1831
rect 4334 1822 4337 1828
rect 1562 1818 2358 1821
rect 2410 1818 4038 1821
rect 802 1808 1318 1811
rect 398 1803 401 1807
rect 397 1802 402 1803
rect 407 1802 408 1807
rect 1422 1803 1425 1807
rect 1421 1802 1426 1803
rect 1431 1802 1432 1807
rect 2446 1803 2449 1807
rect 2445 1802 2450 1803
rect 2455 1802 2456 1807
rect 3478 1803 3481 1807
rect 3477 1802 3482 1803
rect 3487 1802 3488 1807
rect 594 1798 1134 1801
rect 2058 1798 2158 1801
rect 4338 1798 4349 1801
rect 4286 1792 4289 1798
rect 18 1788 854 1791
rect 2226 1788 3702 1791
rect 4346 1788 4349 1791
rect 722 1778 1878 1781
rect 1994 1778 2510 1781
rect 2514 1778 2790 1781
rect 4258 1778 4342 1781
rect 826 1768 1286 1771
rect 1546 1768 2086 1771
rect 2266 1768 3526 1771
rect 1674 1758 2062 1761
rect 2466 1758 3214 1761
rect 3634 1758 3654 1761
rect 3922 1758 4166 1761
rect 1386 1748 1510 1751
rect 2050 1748 2190 1751
rect 2210 1748 3414 1751
rect 4058 1748 4254 1751
rect 170 1738 1230 1741
rect 1722 1738 2014 1741
rect 2018 1738 2046 1741
rect 2066 1738 3758 1741
rect 914 1728 1302 1731
rect 1978 1728 2254 1731
rect 3138 1728 4030 1731
rect 4178 1728 4302 1731
rect 610 1718 1142 1721
rect 1242 1718 1382 1721
rect 1578 1718 1798 1721
rect 1890 1718 2102 1721
rect 3114 1718 4033 1721
rect 1530 1708 1790 1711
rect 1962 1708 2205 1711
rect 3090 1708 3790 1711
rect 4030 1711 4033 1718
rect 4030 1708 4246 1711
rect 902 1703 905 1707
rect 901 1702 906 1703
rect 911 1702 912 1707
rect 1934 1703 1937 1707
rect 1933 1702 1938 1703
rect 1943 1702 1944 1707
rect 2958 1703 2961 1707
rect 2957 1702 2962 1703
rect 2967 1702 2968 1707
rect 3982 1703 3985 1707
rect 3981 1702 3986 1703
rect 3991 1702 3992 1707
rect 2258 1698 2654 1701
rect 3394 1698 3830 1701
rect 4210 1698 4230 1701
rect 722 1688 974 1691
rect 1282 1688 1382 1691
rect 1802 1688 2734 1691
rect 2754 1688 4142 1691
rect 554 1678 2206 1681
rect 2226 1678 3446 1681
rect 3490 1678 3950 1681
rect 158 1671 161 1678
rect 158 1668 1134 1671
rect 1170 1668 1446 1671
rect 1610 1668 1806 1671
rect 1930 1668 2006 1671
rect 2018 1668 3694 1671
rect 3698 1668 3750 1671
rect 1370 1658 2590 1661
rect 794 1648 1078 1651
rect 1122 1648 1510 1651
rect 1682 1648 2169 1651
rect 2386 1648 3158 1651
rect 3170 1648 3246 1651
rect 3306 1648 4118 1651
rect 1922 1638 2006 1641
rect 2166 1641 2169 1648
rect 2166 1638 2870 1641
rect 2882 1638 3470 1641
rect 818 1628 1550 1631
rect 1810 1628 1974 1631
rect 2834 1628 3182 1631
rect 3186 1628 3214 1631
rect 1338 1618 1870 1621
rect 2386 1618 3094 1621
rect 3106 1618 3926 1621
rect 1650 1608 2078 1611
rect 398 1603 401 1607
rect 397 1602 402 1603
rect 407 1602 408 1607
rect 1422 1603 1425 1607
rect 1421 1602 1426 1603
rect 1431 1602 1432 1607
rect 2446 1603 2449 1607
rect 2445 1602 2450 1603
rect 2455 1602 2456 1607
rect 3478 1603 3481 1607
rect 3477 1602 3482 1603
rect 3487 1602 3488 1607
rect 1442 1598 1966 1601
rect 1970 1588 1997 1591
rect 2794 1588 3310 1591
rect 1890 1578 2982 1581
rect 3170 1578 3934 1581
rect 986 1568 1366 1571
rect 1642 1568 1825 1571
rect 1874 1568 2142 1571
rect 2202 1568 3950 1571
rect 1466 1558 1654 1561
rect 1746 1558 1814 1561
rect 1822 1561 1825 1568
rect 4162 1568 4190 1571
rect 1822 1558 1974 1561
rect 2010 1558 3102 1561
rect 3322 1558 3398 1561
rect 3586 1558 3830 1561
rect 818 1548 894 1551
rect 1130 1548 1478 1551
rect 1514 1548 2326 1551
rect 2330 1548 2598 1551
rect 3210 1548 3366 1551
rect 3370 1548 3542 1551
rect 3546 1548 3830 1551
rect 1378 1538 2102 1541
rect 2106 1538 2566 1541
rect 2578 1538 2622 1541
rect 2826 1538 3238 1541
rect 3354 1538 3497 1541
rect 3506 1538 4174 1541
rect 882 1528 1550 1531
rect 1610 1528 1758 1531
rect 1930 1528 2782 1531
rect 2786 1528 3150 1531
rect 3178 1528 3334 1531
rect 3338 1528 3374 1531
rect 3494 1531 3497 1538
rect 3494 1528 3526 1531
rect 3698 1528 3766 1531
rect 594 1518 1518 1521
rect 1682 1518 1886 1521
rect 1918 1518 2830 1521
rect 2858 1518 4046 1521
rect 1918 1511 1921 1518
rect 1098 1508 1921 1511
rect 2426 1508 2942 1511
rect 2986 1508 3118 1511
rect 3122 1508 3470 1511
rect 902 1503 905 1507
rect 901 1502 906 1503
rect 911 1502 912 1507
rect 1934 1503 1937 1507
rect 1933 1502 1938 1503
rect 1943 1502 1944 1507
rect 2958 1503 2961 1507
rect 2957 1502 2962 1503
rect 2967 1502 2968 1507
rect 3982 1503 3985 1507
rect 3981 1502 3986 1503
rect 3991 1502 3992 1507
rect 1562 1498 1894 1501
rect 890 1488 2302 1491
rect 2874 1488 3542 1491
rect 602 1478 838 1481
rect 1106 1478 1494 1481
rect 1690 1478 1894 1481
rect 1914 1478 2342 1481
rect 3226 1478 3310 1481
rect 178 1468 510 1471
rect 514 1468 646 1471
rect 762 1468 1030 1471
rect 1698 1468 1726 1471
rect 1762 1468 2398 1471
rect 2418 1468 2726 1471
rect 2826 1468 3294 1471
rect 3298 1468 3422 1471
rect 4234 1468 4262 1471
rect 202 1458 606 1461
rect 1506 1458 2894 1461
rect 3018 1458 3382 1461
rect 1586 1448 1590 1451
rect 1642 1448 1798 1451
rect 2018 1448 3110 1451
rect 3330 1448 3374 1451
rect 82 1438 710 1441
rect 1682 1438 1913 1441
rect 1930 1438 2886 1441
rect 4002 1438 4094 1441
rect 1910 1432 1913 1438
rect 1762 1428 1838 1431
rect 2434 1428 2846 1431
rect 1570 1418 1926 1421
rect 2266 1418 3622 1421
rect 1650 1408 1654 1411
rect 1658 1408 2429 1411
rect 398 1403 401 1407
rect 397 1402 402 1403
rect 407 1402 408 1407
rect 1422 1403 1425 1407
rect 1421 1402 1426 1403
rect 1431 1402 1432 1407
rect 2446 1403 2449 1407
rect 2445 1402 2450 1403
rect 2455 1402 2456 1407
rect 3478 1403 3481 1407
rect 3477 1402 3482 1403
rect 3487 1402 3488 1407
rect 1730 1398 1822 1401
rect 1498 1388 1998 1391
rect 2346 1388 2526 1391
rect 842 1378 1342 1381
rect 1530 1378 1942 1381
rect 1946 1378 2062 1381
rect 2066 1378 2110 1381
rect 2482 1378 4014 1381
rect 1330 1368 1486 1371
rect 1874 1368 4046 1371
rect 770 1358 918 1361
rect 922 1358 1214 1361
rect 1466 1358 1614 1361
rect 1642 1358 1878 1361
rect 2106 1358 4126 1361
rect 114 1348 966 1351
rect 1282 1348 1374 1351
rect 1418 1348 1574 1351
rect 1602 1348 1670 1351
rect 2010 1348 2070 1351
rect 2074 1348 2326 1351
rect 3546 1348 3646 1351
rect 530 1338 926 1341
rect 1266 1338 1350 1341
rect 1514 1338 1517 1341
rect 1554 1338 2134 1341
rect 2838 1338 3342 1341
rect 3362 1338 3670 1341
rect 250 1328 750 1331
rect 1234 1328 1486 1331
rect 1578 1328 1718 1331
rect 1726 1328 1734 1331
rect 514 1318 918 1321
rect 1010 1318 1310 1321
rect 1394 1318 1526 1321
rect 1534 1318 1549 1321
rect 1534 1311 1537 1318
rect 1726 1321 1729 1328
rect 1618 1318 1729 1321
rect 1766 1321 1769 1328
rect 2838 1331 2841 1338
rect 1794 1328 2841 1331
rect 2850 1328 4150 1331
rect 1738 1318 1769 1321
rect 1842 1318 2798 1321
rect 3290 1318 3622 1321
rect 1346 1308 1537 1311
rect 1554 1308 1638 1311
rect 1722 1308 1789 1311
rect 902 1303 905 1307
rect 901 1302 906 1303
rect 911 1302 912 1307
rect 1210 1298 1542 1301
rect 1638 1301 1641 1308
rect 1826 1308 1910 1311
rect 2018 1308 2126 1311
rect 2434 1308 2638 1311
rect 3314 1308 3326 1311
rect 3330 1308 3502 1311
rect 1934 1303 1937 1307
rect 1933 1302 1938 1303
rect 1943 1302 1944 1307
rect 2958 1303 2961 1307
rect 2957 1302 2962 1303
rect 2967 1302 2968 1307
rect 3982 1303 3985 1307
rect 3981 1302 3986 1303
rect 3991 1302 3992 1307
rect 1638 1298 1837 1301
rect 2022 1298 2870 1301
rect 2874 1298 2926 1301
rect 2978 1298 3422 1301
rect 674 1288 1102 1291
rect 2022 1291 2025 1298
rect 1386 1288 2025 1291
rect 2306 1288 2414 1291
rect 2530 1288 3870 1291
rect 4222 1282 4225 1288
rect 26 1278 678 1281
rect 682 1278 1374 1281
rect 1386 1278 1590 1281
rect 1610 1278 1622 1281
rect 1746 1278 1886 1281
rect 2042 1278 2941 1281
rect 3698 1278 3878 1281
rect 930 1268 1894 1271
rect 2202 1268 2534 1271
rect 2738 1268 2774 1271
rect 3258 1268 3438 1271
rect 3442 1268 3774 1271
rect 4018 1268 4077 1271
rect 506 1258 534 1261
rect 1298 1258 1414 1261
rect 1474 1258 1798 1261
rect 1802 1258 2142 1261
rect 2290 1258 3254 1261
rect 3626 1258 3758 1261
rect 1330 1248 1533 1251
rect 1546 1248 1750 1251
rect 1762 1248 2510 1251
rect 2946 1248 4054 1251
rect 18 1238 926 1241
rect 1058 1238 1982 1241
rect 1986 1238 2102 1241
rect 2202 1238 2710 1241
rect 2714 1238 3246 1241
rect 3370 1238 4286 1241
rect 1498 1228 1534 1231
rect 1554 1228 1766 1231
rect 1826 1228 3070 1231
rect 1362 1218 1750 1221
rect 1786 1218 1901 1221
rect 2002 1218 2318 1221
rect 2430 1218 2902 1221
rect 2906 1218 3198 1221
rect 3242 1218 3726 1221
rect 810 1208 1078 1211
rect 1442 1208 2270 1211
rect 2430 1211 2433 1218
rect 2274 1208 2433 1211
rect 2842 1208 3197 1211
rect 398 1203 401 1207
rect 397 1202 402 1203
rect 407 1202 408 1207
rect 1422 1203 1425 1207
rect 1421 1202 1426 1203
rect 1431 1202 1432 1207
rect 2446 1203 2449 1207
rect 2445 1202 2450 1203
rect 2455 1202 2456 1207
rect 3478 1203 3481 1207
rect 3477 1202 3482 1203
rect 3487 1202 3488 1207
rect 930 1198 1382 1201
rect 1538 1198 2238 1201
rect 698 1188 1118 1191
rect 1394 1188 1822 1191
rect 2122 1188 3062 1191
rect 3450 1188 3622 1191
rect 26 1178 758 1181
rect 762 1178 1102 1181
rect 1106 1178 1182 1181
rect 1578 1178 1613 1181
rect 1634 1178 1725 1181
rect 1922 1178 2222 1181
rect 2242 1178 3710 1181
rect 1234 1168 2350 1171
rect 3562 1168 3782 1171
rect 690 1158 926 1161
rect 754 1148 934 1151
rect 1070 1151 1073 1158
rect 2194 1158 2566 1161
rect 2570 1158 3062 1161
rect 4286 1161 4289 1168
rect 3210 1158 4289 1161
rect 3102 1152 3105 1158
rect 1070 1148 1198 1151
rect 1378 1148 2790 1151
rect 3490 1148 3998 1151
rect 1210 1138 2189 1141
rect 2202 1138 3110 1141
rect 3114 1138 3254 1141
rect 658 1128 974 1131
rect 1234 1128 1238 1131
rect 1282 1128 1398 1131
rect 1562 1128 1581 1131
rect 1626 1128 1998 1131
rect 2026 1128 2638 1131
rect 2658 1128 2822 1131
rect 3018 1128 3053 1131
rect 3150 1128 3230 1131
rect 3762 1128 3886 1131
rect 1534 1122 1537 1127
rect 3150 1122 3153 1128
rect 1706 1118 2702 1121
rect 2738 1118 3006 1121
rect 4306 1118 4334 1121
rect 1210 1108 1622 1111
rect 3002 1108 3958 1111
rect 4306 1108 4350 1111
rect 902 1103 905 1107
rect 901 1102 906 1103
rect 911 1102 912 1107
rect 1934 1103 1937 1107
rect 1933 1102 1938 1103
rect 1943 1102 1944 1107
rect 2958 1103 2961 1107
rect 2957 1102 2962 1103
rect 2967 1102 2968 1107
rect 3982 1103 3985 1107
rect 3981 1102 3986 1103
rect 3991 1102 3992 1107
rect 1274 1098 1774 1101
rect 1050 1088 1534 1091
rect 1666 1088 1774 1091
rect 1826 1088 2198 1091
rect 2890 1088 2982 1091
rect 3018 1088 4222 1091
rect 938 1078 1262 1081
rect 1354 1078 1478 1081
rect 1482 1078 1542 1081
rect 1566 1081 1569 1088
rect 4290 1088 4358 1091
rect 1566 1078 1854 1081
rect 1866 1078 2126 1081
rect 2362 1078 3086 1081
rect 3114 1078 3446 1081
rect 170 1068 702 1071
rect 1082 1068 1437 1071
rect 982 1061 985 1068
rect 1626 1068 1702 1071
rect 1770 1068 3734 1071
rect 982 1058 1302 1061
rect 1314 1058 1710 1061
rect 1858 1058 2550 1061
rect 2778 1058 3262 1061
rect 3594 1058 3710 1061
rect 3962 1058 4142 1061
rect 778 1048 1150 1051
rect 1474 1048 2270 1051
rect 2282 1048 2366 1051
rect 2522 1048 2942 1051
rect 2946 1048 3334 1051
rect 3474 1048 3830 1051
rect 4170 1048 4246 1051
rect 1658 1038 2030 1041
rect 2146 1038 2998 1041
rect 3090 1038 3526 1041
rect 4178 1038 4238 1041
rect 1466 1028 1638 1031
rect 2410 1028 3814 1031
rect 4270 1022 4273 1027
rect 1042 1018 2190 1021
rect 2342 1018 3062 1021
rect 3066 1018 3198 1021
rect 3462 1018 4222 1021
rect 2342 1011 2345 1018
rect 1714 1008 2345 1011
rect 2754 1008 2878 1011
rect 3462 1011 3465 1018
rect 3002 1008 3465 1011
rect 4194 1008 4222 1011
rect 398 1003 401 1007
rect 397 1002 402 1003
rect 407 1002 408 1007
rect 1422 1003 1425 1007
rect 1421 1002 1426 1003
rect 1431 1002 1432 1007
rect 2446 1003 2449 1007
rect 2445 1002 2450 1003
rect 2455 1002 2456 1007
rect 3478 1003 3481 1007
rect 3477 1002 3482 1003
rect 3487 1002 3488 1007
rect 1490 988 1510 991
rect 1522 988 3150 991
rect 1042 978 1686 981
rect 1690 978 2541 981
rect 2562 978 3126 981
rect 522 968 1254 971
rect 1258 968 1501 971
rect 1514 968 1854 971
rect 1874 968 1990 971
rect 2026 968 4214 971
rect 666 958 1222 961
rect 1754 958 2054 961
rect 2250 958 2510 961
rect 2634 958 3134 961
rect 1138 948 1150 951
rect 1210 948 1262 951
rect 1506 948 2046 951
rect 2054 951 2057 958
rect 2054 948 4246 951
rect 1234 938 2502 941
rect 2506 938 3070 941
rect 3074 938 3622 941
rect 3762 938 3814 941
rect 1338 928 1654 931
rect 1658 928 2118 931
rect 3306 928 3414 931
rect 3594 928 3766 931
rect 3770 928 3998 931
rect 1330 918 1550 921
rect 1554 918 1870 921
rect 1890 918 3310 921
rect 3354 918 3422 921
rect 1538 908 1542 911
rect 1562 908 1869 911
rect 902 903 905 907
rect 901 902 906 903
rect 911 902 912 907
rect 1934 903 1937 907
rect 1933 902 1938 903
rect 1943 902 1944 907
rect 2958 903 2961 907
rect 2957 902 2962 903
rect 2967 902 2968 907
rect 3982 903 3985 907
rect 3981 902 3986 903
rect 3991 902 3992 907
rect 1026 898 1398 901
rect 2394 898 2886 901
rect 3122 898 3318 901
rect 1402 888 1726 891
rect 1874 888 3086 891
rect 3106 888 3958 891
rect 1146 878 1686 881
rect 1730 878 1830 881
rect 2226 878 2526 881
rect 2586 878 2670 881
rect 2890 878 4110 881
rect 4146 878 4206 881
rect 170 868 814 871
rect 1402 868 1454 871
rect 1658 868 1726 871
rect 1766 868 2318 871
rect 2322 868 2774 871
rect 2946 868 3926 871
rect 762 858 1278 861
rect 1454 861 1457 868
rect 1766 861 1769 868
rect 1454 858 1769 861
rect 2178 858 2934 861
rect 3194 858 3398 861
rect 3402 858 3686 861
rect 826 848 974 851
rect 1458 848 1942 851
rect 2626 848 4310 851
rect 1354 838 1582 841
rect 1906 838 1974 841
rect 2290 838 2766 841
rect 3186 838 3902 841
rect 1674 828 2670 831
rect 2898 828 3198 831
rect 1386 818 1854 821
rect 1858 818 2918 821
rect 2978 818 3502 821
rect 1498 808 1862 811
rect 1874 808 1910 811
rect 2546 808 2566 811
rect 2570 808 2710 811
rect 2714 808 3078 811
rect 398 803 401 807
rect 397 802 402 803
rect 407 802 408 807
rect 1422 803 1425 807
rect 1421 802 1426 803
rect 1431 802 1432 807
rect 2446 803 2449 807
rect 2445 802 2450 803
rect 2455 802 2456 807
rect 3478 803 3481 807
rect 3477 802 3482 803
rect 3487 802 3488 807
rect 1522 798 1590 801
rect 1698 798 1702 801
rect 1554 788 1798 791
rect 1802 788 3134 791
rect 3306 788 3566 791
rect 1434 778 1990 781
rect 2066 778 4206 781
rect 4210 778 4254 781
rect 1426 768 2086 771
rect 2402 768 2662 771
rect 2778 768 3366 771
rect 1722 758 2061 761
rect 2074 758 2654 761
rect 2730 758 4102 761
rect 1370 748 1705 751
rect 2042 748 3934 751
rect 4058 748 4093 751
rect 1702 742 1705 748
rect 170 738 1134 741
rect 2034 738 2486 741
rect 2490 738 2678 741
rect 3114 738 3806 741
rect 1618 728 1662 731
rect 2514 728 2518 731
rect 2602 728 2694 731
rect 3642 728 4006 731
rect 1698 718 2358 721
rect 2530 718 2718 721
rect 2882 718 3510 721
rect 1466 708 1582 711
rect 1650 708 1902 711
rect 2410 708 2886 711
rect 3162 708 3422 711
rect 902 703 905 707
rect 901 702 906 703
rect 911 702 912 707
rect 1934 703 1937 707
rect 1933 702 1938 703
rect 1943 702 1944 707
rect 2958 703 2961 707
rect 2957 702 2962 703
rect 2967 702 2968 707
rect 3982 703 3985 707
rect 3981 702 3986 703
rect 3991 702 3992 707
rect 1466 698 1846 701
rect 3266 698 3430 701
rect 138 688 918 691
rect 1778 688 3302 691
rect 3394 688 3710 691
rect 1314 678 1614 681
rect 3234 678 3502 681
rect 394 668 942 671
rect 2110 671 2113 678
rect 1258 668 1489 671
rect 2110 668 2206 671
rect 2322 668 3246 671
rect 3546 668 3878 671
rect 1486 662 1489 668
rect 4078 662 4081 668
rect 1490 658 2590 661
rect 2626 658 2726 661
rect 3370 658 3702 661
rect 1410 648 2414 651
rect 2426 648 2926 651
rect 2930 648 3006 651
rect 3202 638 4302 641
rect 1906 628 2894 631
rect 1562 618 2918 621
rect 398 603 401 607
rect 397 602 402 603
rect 407 602 408 607
rect 1422 603 1425 607
rect 1421 602 1426 603
rect 1431 602 1432 607
rect 2446 603 2449 607
rect 2445 602 2450 603
rect 2455 602 2456 607
rect 3478 603 3481 607
rect 3477 602 3482 603
rect 3487 602 3488 607
rect 1602 598 2422 601
rect 2682 588 3238 591
rect 1666 578 1974 581
rect 2178 578 3902 581
rect 1462 568 1854 571
rect 1986 568 4078 571
rect 1462 562 1465 568
rect 2210 558 2614 561
rect 2618 558 2774 561
rect 3218 558 4070 561
rect 1418 548 1982 551
rect 2834 548 3937 551
rect 3934 542 3937 548
rect 2018 528 3246 531
rect 3298 528 4110 531
rect 2002 518 3902 521
rect 2266 508 2534 511
rect 3002 508 3230 511
rect 3234 508 3726 511
rect 902 503 905 507
rect 901 502 906 503
rect 911 502 912 507
rect 1934 503 1937 507
rect 1933 502 1938 503
rect 1943 502 1944 507
rect 2958 503 2961 507
rect 2957 502 2962 503
rect 2967 502 2968 507
rect 3982 503 3985 507
rect 3981 502 3986 503
rect 3991 502 3992 507
rect 2954 488 3182 491
rect 1222 481 1225 488
rect 1222 478 1294 481
rect 1450 478 2046 481
rect 2114 478 2678 481
rect 3098 478 3118 481
rect 4346 478 4349 481
rect 1762 468 3998 471
rect 1778 458 3310 461
rect 2322 448 2518 451
rect 2526 448 2534 451
rect 2538 448 2774 451
rect 3010 448 3094 451
rect 3898 448 4326 451
rect 2394 438 2926 441
rect 3122 438 3670 441
rect 1202 428 1542 431
rect 1546 428 2462 431
rect 3998 422 4001 427
rect 2546 408 3326 411
rect 398 403 401 407
rect 397 402 402 403
rect 407 402 408 407
rect 1422 403 1425 407
rect 1421 402 1426 403
rect 1431 402 1432 407
rect 2446 403 2449 407
rect 2445 402 2450 403
rect 2455 402 2456 407
rect 3478 403 3481 407
rect 3477 402 3482 403
rect 3487 402 3488 407
rect 778 398 1230 401
rect 1746 398 2398 401
rect 2522 398 3053 401
rect 3058 398 3262 401
rect 1490 388 2022 391
rect 2498 388 4078 391
rect 2338 378 2534 381
rect 2538 378 3230 381
rect 1802 368 2054 371
rect 3858 368 3942 371
rect 1522 358 3254 361
rect 3706 358 3910 361
rect 3954 358 4289 361
rect 4286 352 4289 358
rect 1314 348 1678 351
rect 1730 348 1942 351
rect 2418 348 2894 351
rect 218 338 1294 341
rect 3718 338 3726 341
rect 3750 341 3753 348
rect 3730 338 3753 341
rect 1834 328 2566 331
rect 2930 328 3886 331
rect 3962 328 4030 331
rect 730 318 1150 321
rect 1354 318 3521 321
rect 3530 318 3726 321
rect 3730 318 3974 321
rect 3518 311 3521 318
rect 3518 308 3886 311
rect 902 303 905 307
rect 901 302 906 303
rect 911 302 912 307
rect 1934 303 1937 307
rect 1933 302 1938 303
rect 1943 302 1944 307
rect 2958 303 2961 307
rect 2957 302 2962 303
rect 2967 302 2968 307
rect 3982 303 3985 307
rect 3981 302 3986 303
rect 3991 302 3992 307
rect 954 298 1270 301
rect 2426 298 2934 301
rect 3410 298 3686 301
rect 2274 288 3137 291
rect 3146 288 4238 291
rect 1786 278 2806 281
rect 3134 281 3137 288
rect 3134 278 3949 281
rect 534 271 537 278
rect 3970 278 4174 281
rect 534 268 918 271
rect 1202 268 1438 271
rect 2386 268 3241 271
rect 4082 268 4085 271
rect 1490 258 2414 261
rect 3238 261 3241 268
rect 3238 258 4070 261
rect 1986 248 2854 251
rect 1482 238 3454 241
rect 3474 238 3902 241
rect 842 228 1229 231
rect 1234 228 1510 231
rect 3426 228 4070 231
rect 2122 218 4062 221
rect 398 203 401 207
rect 397 202 402 203
rect 407 202 408 207
rect 1422 203 1425 207
rect 1421 202 1426 203
rect 1431 202 1432 207
rect 2446 203 2449 207
rect 2445 202 2450 203
rect 2455 202 2456 207
rect 3478 203 3481 207
rect 3477 202 3482 203
rect 3487 202 3488 207
rect 1610 198 2262 201
rect 1314 188 2286 191
rect 2330 188 4206 191
rect 2218 178 2534 181
rect 2538 178 3574 181
rect 3578 178 3638 181
rect 498 168 1214 171
rect 2010 168 3454 171
rect 698 158 1118 161
rect 1282 158 2126 161
rect 4242 158 4294 161
rect 4370 158 4381 161
rect 218 148 990 151
rect 1154 148 1254 151
rect 1406 148 1606 151
rect 1930 148 2078 151
rect 2226 148 2702 151
rect 2706 148 3830 151
rect 4306 148 4365 151
rect 1406 142 1409 148
rect 1122 138 1310 141
rect 1554 138 1638 141
rect 1714 138 2422 141
rect 4302 132 4305 138
rect 1090 128 1262 131
rect 1378 128 2094 131
rect 2498 128 2566 131
rect 2570 128 2662 131
rect 2698 128 3182 131
rect 4322 128 4326 131
rect 1394 118 3350 121
rect 4178 108 4221 111
rect 902 103 905 107
rect 901 102 906 103
rect 911 102 912 107
rect 1934 103 1937 107
rect 1933 102 1938 103
rect 1943 102 1944 107
rect 2958 103 2961 107
rect 2957 102 2962 103
rect 2967 102 2968 107
rect 3982 103 3985 107
rect 3981 102 3986 103
rect 3991 102 3992 107
rect 4130 98 4150 101
rect 162 88 1342 91
rect 1594 88 2974 91
rect 4202 88 4205 91
rect 4142 82 4145 87
rect 1258 78 1438 81
rect 1506 78 2718 81
rect 1102 71 1105 78
rect 1102 68 1238 71
rect 1242 68 2054 71
rect 2610 68 3174 71
rect 3594 68 3686 71
rect 4322 68 4333 71
rect 554 58 1382 61
rect 1570 58 3726 61
rect 4162 38 4174 41
rect 1338 28 2174 31
rect 1426 18 2086 21
rect 398 3 401 7
rect 397 2 402 3
rect 407 2 408 7
rect 1422 3 1425 7
rect 1421 2 1426 3
rect 1431 2 1432 7
rect 2446 3 2449 7
rect 2445 2 2450 3
rect 2455 2 2456 7
rect 3478 3 3481 7
rect 3477 2 3482 3
rect 3487 2 3488 7
<< m6contact >>
rect 896 3103 898 3107
rect 898 3103 901 3107
rect 906 3103 909 3107
rect 909 3103 911 3107
rect 896 3102 901 3103
rect 906 3102 911 3103
rect 1928 3103 1930 3107
rect 1930 3103 1933 3107
rect 1938 3103 1941 3107
rect 1941 3103 1943 3107
rect 1928 3102 1933 3103
rect 1938 3102 1943 3103
rect 2952 3103 2954 3107
rect 2954 3103 2957 3107
rect 2962 3103 2965 3107
rect 2965 3103 2967 3107
rect 2952 3102 2957 3103
rect 2962 3102 2967 3103
rect 3976 3103 3978 3107
rect 3978 3103 3981 3107
rect 3986 3103 3989 3107
rect 3989 3103 3991 3107
rect 3976 3102 3981 3103
rect 3986 3102 3991 3103
rect 4301 3067 4306 3072
rect 4253 3047 4258 3052
rect 4269 3037 4274 3042
rect 392 3003 394 3007
rect 394 3003 397 3007
rect 402 3003 405 3007
rect 405 3003 407 3007
rect 392 3002 397 3003
rect 402 3002 407 3003
rect 1416 3003 1418 3007
rect 1418 3003 1421 3007
rect 1426 3003 1429 3007
rect 1429 3003 1431 3007
rect 1416 3002 1421 3003
rect 1426 3002 1431 3003
rect 2440 3003 2442 3007
rect 2442 3003 2445 3007
rect 2450 3003 2453 3007
rect 2453 3003 2455 3007
rect 2440 3002 2445 3003
rect 2450 3002 2455 3003
rect 3472 3003 3474 3007
rect 3474 3003 3477 3007
rect 3482 3003 3485 3007
rect 3485 3003 3487 3007
rect 3472 3002 3477 3003
rect 3482 3002 3487 3003
rect 896 2903 898 2907
rect 898 2903 901 2907
rect 906 2903 909 2907
rect 909 2903 911 2907
rect 896 2902 901 2903
rect 906 2902 911 2903
rect 1928 2903 1930 2907
rect 1930 2903 1933 2907
rect 1938 2903 1941 2907
rect 1941 2903 1943 2907
rect 1928 2902 1933 2903
rect 1938 2902 1943 2903
rect 2952 2903 2954 2907
rect 2954 2903 2957 2907
rect 2962 2903 2965 2907
rect 2965 2903 2967 2907
rect 2952 2902 2957 2903
rect 2962 2902 2967 2903
rect 3976 2903 3978 2907
rect 3978 2903 3981 2907
rect 3986 2903 3989 2907
rect 3989 2903 3991 2907
rect 3976 2902 3981 2903
rect 3986 2902 3991 2903
rect 392 2803 394 2807
rect 394 2803 397 2807
rect 402 2803 405 2807
rect 405 2803 407 2807
rect 392 2802 397 2803
rect 402 2802 407 2803
rect 1416 2803 1418 2807
rect 1418 2803 1421 2807
rect 1426 2803 1429 2807
rect 1429 2803 1431 2807
rect 1416 2802 1421 2803
rect 1426 2802 1431 2803
rect 2440 2803 2442 2807
rect 2442 2803 2445 2807
rect 2450 2803 2453 2807
rect 2453 2803 2455 2807
rect 2440 2802 2445 2803
rect 2450 2802 2455 2803
rect 3472 2803 3474 2807
rect 3474 2803 3477 2807
rect 3482 2803 3485 2807
rect 3485 2803 3487 2807
rect 3472 2802 3477 2803
rect 3482 2802 3487 2803
rect 4125 2767 4130 2772
rect 3197 2757 3202 2762
rect 4349 2747 4354 2752
rect 4317 2737 4322 2742
rect 896 2703 898 2707
rect 898 2703 901 2707
rect 906 2703 909 2707
rect 909 2703 911 2707
rect 896 2702 901 2703
rect 906 2702 911 2703
rect 1928 2703 1930 2707
rect 1930 2703 1933 2707
rect 1938 2703 1941 2707
rect 1941 2703 1943 2707
rect 1928 2702 1933 2703
rect 1938 2702 1943 2703
rect 2952 2703 2954 2707
rect 2954 2703 2957 2707
rect 2962 2703 2965 2707
rect 2965 2703 2967 2707
rect 2952 2702 2957 2703
rect 2962 2702 2967 2703
rect 3976 2703 3978 2707
rect 3978 2703 3981 2707
rect 3986 2703 3989 2707
rect 3989 2703 3991 2707
rect 3976 2702 3981 2703
rect 3986 2702 3991 2703
rect 4301 2647 4306 2652
rect 392 2603 394 2607
rect 394 2603 397 2607
rect 402 2603 405 2607
rect 405 2603 407 2607
rect 392 2602 397 2603
rect 402 2602 407 2603
rect 1416 2603 1418 2607
rect 1418 2603 1421 2607
rect 1426 2603 1429 2607
rect 1429 2603 1431 2607
rect 1416 2602 1421 2603
rect 1426 2602 1431 2603
rect 2440 2603 2442 2607
rect 2442 2603 2445 2607
rect 2450 2603 2453 2607
rect 2453 2603 2455 2607
rect 2440 2602 2445 2603
rect 2450 2602 2455 2603
rect 3472 2603 3474 2607
rect 3474 2603 3477 2607
rect 3482 2603 3485 2607
rect 3485 2603 3487 2607
rect 3472 2602 3477 2603
rect 3482 2602 3487 2603
rect 896 2503 898 2507
rect 898 2503 901 2507
rect 906 2503 909 2507
rect 909 2503 911 2507
rect 896 2502 901 2503
rect 906 2502 911 2503
rect 1928 2503 1930 2507
rect 1930 2503 1933 2507
rect 1938 2503 1941 2507
rect 1941 2503 1943 2507
rect 1928 2502 1933 2503
rect 1938 2502 1943 2503
rect 2952 2503 2954 2507
rect 2954 2503 2957 2507
rect 2962 2503 2965 2507
rect 2965 2503 2967 2507
rect 2952 2502 2957 2503
rect 2962 2502 2967 2503
rect 3976 2503 3978 2507
rect 3978 2503 3981 2507
rect 3986 2503 3989 2507
rect 3989 2503 3991 2507
rect 3976 2502 3981 2503
rect 3986 2502 3991 2503
rect 2941 2497 2946 2502
rect 2941 2467 2946 2472
rect 3101 2467 3106 2472
rect 4365 2437 4370 2442
rect 1997 2427 2002 2432
rect 392 2403 394 2407
rect 394 2403 397 2407
rect 402 2403 405 2407
rect 405 2403 407 2407
rect 392 2402 397 2403
rect 402 2402 407 2403
rect 1416 2403 1418 2407
rect 1418 2403 1421 2407
rect 1426 2403 1429 2407
rect 1429 2403 1431 2407
rect 1416 2402 1421 2403
rect 1426 2402 1431 2403
rect 2440 2403 2442 2407
rect 2442 2403 2445 2407
rect 2450 2403 2453 2407
rect 2453 2403 2455 2407
rect 2440 2402 2445 2403
rect 2450 2402 2455 2403
rect 3472 2403 3474 2407
rect 3474 2403 3477 2407
rect 3482 2403 3485 2407
rect 3485 2403 3487 2407
rect 3472 2402 3477 2403
rect 3482 2402 3487 2403
rect 4381 2357 4386 2362
rect 1869 2347 1874 2352
rect 1997 2347 2002 2352
rect 4301 2347 4306 2352
rect 1869 2317 1874 2322
rect 896 2303 898 2307
rect 898 2303 901 2307
rect 906 2303 909 2307
rect 909 2303 911 2307
rect 896 2302 901 2303
rect 906 2302 911 2303
rect 1928 2303 1930 2307
rect 1930 2303 1933 2307
rect 1938 2303 1941 2307
rect 1941 2303 1943 2307
rect 1928 2302 1933 2303
rect 1938 2302 1943 2303
rect 2952 2303 2954 2307
rect 2954 2303 2957 2307
rect 2962 2303 2965 2307
rect 2965 2303 2967 2307
rect 2952 2302 2957 2303
rect 2962 2302 2967 2303
rect 3976 2303 3978 2307
rect 3978 2303 3981 2307
rect 3986 2303 3989 2307
rect 3989 2303 3991 2307
rect 3976 2302 3981 2303
rect 3986 2302 3991 2303
rect 392 2203 394 2207
rect 394 2203 397 2207
rect 402 2203 405 2207
rect 405 2203 407 2207
rect 392 2202 397 2203
rect 402 2202 407 2203
rect 1416 2203 1418 2207
rect 1418 2203 1421 2207
rect 1426 2203 1429 2207
rect 1429 2203 1431 2207
rect 1416 2202 1421 2203
rect 1426 2202 1431 2203
rect 2440 2203 2442 2207
rect 2442 2203 2445 2207
rect 2450 2203 2453 2207
rect 2453 2203 2455 2207
rect 2440 2202 2445 2203
rect 2450 2202 2455 2203
rect 3472 2203 3474 2207
rect 3474 2203 3477 2207
rect 3482 2203 3485 2207
rect 3485 2203 3487 2207
rect 3472 2202 3477 2203
rect 3482 2202 3487 2203
rect 3277 2187 3282 2192
rect 4077 2147 4082 2152
rect 4093 2147 4098 2152
rect 896 2103 898 2107
rect 898 2103 901 2107
rect 906 2103 909 2107
rect 909 2103 911 2107
rect 896 2102 901 2103
rect 906 2102 911 2103
rect 1928 2103 1930 2107
rect 1930 2103 1933 2107
rect 1938 2103 1941 2107
rect 1941 2103 1943 2107
rect 1928 2102 1933 2103
rect 1938 2102 1943 2103
rect 2952 2103 2954 2107
rect 2954 2103 2957 2107
rect 2962 2103 2965 2107
rect 2965 2103 2967 2107
rect 2952 2102 2957 2103
rect 2962 2102 2967 2103
rect 3976 2103 3978 2107
rect 3978 2103 3981 2107
rect 3986 2103 3989 2107
rect 3989 2103 3991 2107
rect 3976 2102 3981 2103
rect 3986 2102 3991 2103
rect 1725 2067 1730 2072
rect 3277 2047 3282 2052
rect 4237 2017 4242 2022
rect 392 2003 394 2007
rect 394 2003 397 2007
rect 402 2003 405 2007
rect 405 2003 407 2007
rect 392 2002 397 2003
rect 402 2002 407 2003
rect 1416 2003 1418 2007
rect 1418 2003 1421 2007
rect 1426 2003 1429 2007
rect 1429 2003 1431 2007
rect 1416 2002 1421 2003
rect 1426 2002 1431 2003
rect 2440 2003 2442 2007
rect 2442 2003 2445 2007
rect 2450 2003 2453 2007
rect 2453 2003 2455 2007
rect 2440 2002 2445 2003
rect 2450 2002 2455 2003
rect 3472 2003 3474 2007
rect 3474 2003 3477 2007
rect 3482 2003 3485 2007
rect 3485 2003 3487 2007
rect 3472 2002 3477 2003
rect 3482 2002 3487 2003
rect 1901 1937 1906 1942
rect 4189 1937 4194 1942
rect 896 1903 898 1907
rect 898 1903 901 1907
rect 906 1903 909 1907
rect 909 1903 911 1907
rect 896 1902 901 1903
rect 906 1902 911 1903
rect 1928 1903 1930 1907
rect 1930 1903 1933 1907
rect 1938 1903 1941 1907
rect 1941 1903 1943 1907
rect 1928 1902 1933 1903
rect 1938 1902 1943 1903
rect 2952 1903 2954 1907
rect 2954 1903 2957 1907
rect 2962 1903 2965 1907
rect 2965 1903 2967 1907
rect 2952 1902 2957 1903
rect 2962 1902 2967 1903
rect 3976 1903 3978 1907
rect 3978 1903 3981 1907
rect 3986 1903 3989 1907
rect 3989 1903 3991 1907
rect 3976 1902 3981 1903
rect 3986 1902 3991 1903
rect 1613 1857 1618 1862
rect 3997 1847 4002 1852
rect 4333 1817 4338 1822
rect 392 1803 394 1807
rect 394 1803 397 1807
rect 402 1803 405 1807
rect 405 1803 407 1807
rect 392 1802 397 1803
rect 402 1802 407 1803
rect 1416 1803 1418 1807
rect 1418 1803 1421 1807
rect 1426 1803 1429 1807
rect 1429 1803 1431 1807
rect 1416 1802 1421 1803
rect 1426 1802 1431 1803
rect 2440 1803 2442 1807
rect 2442 1803 2445 1807
rect 2450 1803 2453 1807
rect 2453 1803 2455 1807
rect 2440 1802 2445 1803
rect 2450 1802 2455 1803
rect 3472 1803 3474 1807
rect 3474 1803 3477 1807
rect 3482 1803 3485 1807
rect 3485 1803 3487 1807
rect 3472 1802 3477 1803
rect 3482 1802 3487 1803
rect 4349 1797 4354 1802
rect 4285 1787 4290 1792
rect 4349 1787 4354 1792
rect 4253 1777 4258 1782
rect 2205 1747 2210 1752
rect 4173 1727 4178 1732
rect 2205 1707 2210 1712
rect 896 1703 898 1707
rect 898 1703 901 1707
rect 906 1703 909 1707
rect 909 1703 911 1707
rect 896 1702 901 1703
rect 906 1702 911 1703
rect 1928 1703 1930 1707
rect 1930 1703 1933 1707
rect 1938 1703 1941 1707
rect 1941 1703 1943 1707
rect 1928 1702 1933 1703
rect 1938 1702 1943 1703
rect 2952 1703 2954 1707
rect 2954 1703 2957 1707
rect 2962 1703 2965 1707
rect 2965 1703 2967 1707
rect 2952 1702 2957 1703
rect 2962 1702 2967 1703
rect 3976 1703 3978 1707
rect 3978 1703 3981 1707
rect 3986 1703 3989 1707
rect 3989 1703 3991 1707
rect 3976 1702 3981 1703
rect 3986 1702 3991 1703
rect 4205 1697 4210 1702
rect 392 1603 394 1607
rect 394 1603 397 1607
rect 402 1603 405 1607
rect 405 1603 407 1607
rect 392 1602 397 1603
rect 402 1602 407 1603
rect 1416 1603 1418 1607
rect 1418 1603 1421 1607
rect 1426 1603 1429 1607
rect 1429 1603 1431 1607
rect 1416 1602 1421 1603
rect 1426 1602 1431 1603
rect 2440 1603 2442 1607
rect 2442 1603 2445 1607
rect 2450 1603 2453 1607
rect 2453 1603 2455 1607
rect 2440 1602 2445 1603
rect 2450 1602 2455 1603
rect 3472 1603 3474 1607
rect 3474 1603 3477 1607
rect 3482 1603 3485 1607
rect 3485 1603 3487 1607
rect 3472 1602 3477 1603
rect 3482 1602 3487 1603
rect 1437 1597 1442 1602
rect 1997 1587 2002 1592
rect 4157 1567 4162 1572
rect 896 1503 898 1507
rect 898 1503 901 1507
rect 906 1503 909 1507
rect 909 1503 911 1507
rect 896 1502 901 1503
rect 906 1502 911 1503
rect 1928 1503 1930 1507
rect 1930 1503 1933 1507
rect 1938 1503 1941 1507
rect 1941 1503 1943 1507
rect 1928 1502 1933 1503
rect 1938 1502 1943 1503
rect 2952 1503 2954 1507
rect 2954 1503 2957 1507
rect 2962 1503 2965 1507
rect 2965 1503 2967 1507
rect 2952 1502 2957 1503
rect 2962 1502 2967 1503
rect 3976 1503 3978 1507
rect 3978 1503 3981 1507
rect 3986 1503 3989 1507
rect 3989 1503 3991 1507
rect 3976 1502 3981 1503
rect 3986 1502 3991 1503
rect 1693 1467 1698 1472
rect 1581 1447 1586 1452
rect 2429 1427 2434 1432
rect 2429 1407 2434 1412
rect 392 1403 394 1407
rect 394 1403 397 1407
rect 402 1403 405 1407
rect 405 1403 407 1407
rect 392 1402 397 1403
rect 402 1402 407 1403
rect 1416 1403 1418 1407
rect 1418 1403 1421 1407
rect 1426 1403 1429 1407
rect 1429 1403 1431 1407
rect 1416 1402 1421 1403
rect 1426 1402 1431 1403
rect 2440 1403 2442 1407
rect 2442 1403 2445 1407
rect 2450 1403 2453 1407
rect 2453 1403 2455 1407
rect 2440 1402 2445 1403
rect 2450 1402 2455 1403
rect 3472 1403 3474 1407
rect 3474 1403 3477 1407
rect 3482 1403 3485 1407
rect 3485 1403 3487 1407
rect 3472 1402 3477 1403
rect 3482 1402 3487 1403
rect 1517 1337 1522 1342
rect 1549 1317 1554 1322
rect 1789 1327 1794 1332
rect 1837 1317 1842 1322
rect 896 1303 898 1307
rect 898 1303 901 1307
rect 906 1303 909 1307
rect 909 1303 911 1307
rect 896 1302 901 1303
rect 906 1302 911 1303
rect 1789 1307 1794 1312
rect 1928 1303 1930 1307
rect 1930 1303 1933 1307
rect 1938 1303 1941 1307
rect 1941 1303 1943 1307
rect 1928 1302 1933 1303
rect 1938 1302 1943 1303
rect 2952 1303 2954 1307
rect 2954 1303 2957 1307
rect 2962 1303 2965 1307
rect 2965 1303 2967 1307
rect 2952 1302 2957 1303
rect 2962 1302 2967 1303
rect 3976 1303 3978 1307
rect 3978 1303 3981 1307
rect 3986 1303 3989 1307
rect 3989 1303 3991 1307
rect 3976 1302 3981 1303
rect 3986 1302 3991 1303
rect 1837 1297 1842 1302
rect 2941 1277 2946 1282
rect 4221 1277 4226 1282
rect 4077 1267 4082 1272
rect 1533 1247 1538 1252
rect 2941 1247 2946 1252
rect 1549 1227 1554 1232
rect 1901 1217 1906 1222
rect 3197 1207 3202 1212
rect 392 1203 394 1207
rect 394 1203 397 1207
rect 402 1203 405 1207
rect 405 1203 407 1207
rect 392 1202 397 1203
rect 402 1202 407 1203
rect 1416 1203 1418 1207
rect 1418 1203 1421 1207
rect 1426 1203 1429 1207
rect 1429 1203 1431 1207
rect 1416 1202 1421 1203
rect 1426 1202 1431 1203
rect 2440 1203 2442 1207
rect 2442 1203 2445 1207
rect 2450 1203 2453 1207
rect 2453 1203 2455 1207
rect 2440 1202 2445 1203
rect 2450 1202 2455 1203
rect 3472 1203 3474 1207
rect 3474 1203 3477 1207
rect 3482 1203 3485 1207
rect 3485 1203 3487 1207
rect 3472 1202 3477 1203
rect 3482 1202 3487 1203
rect 1533 1197 1538 1202
rect 1613 1177 1618 1182
rect 1725 1177 1730 1182
rect 2189 1157 2194 1162
rect 3101 1147 3106 1152
rect 2189 1137 2194 1142
rect 1229 1127 1234 1132
rect 1533 1127 1538 1132
rect 1581 1127 1586 1132
rect 3053 1127 3058 1132
rect 4301 1117 4306 1122
rect 4301 1107 4306 1112
rect 896 1103 898 1107
rect 898 1103 901 1107
rect 906 1103 909 1107
rect 909 1103 911 1107
rect 896 1102 901 1103
rect 906 1102 911 1103
rect 1928 1103 1930 1107
rect 1930 1103 1933 1107
rect 1938 1103 1941 1107
rect 1941 1103 1943 1107
rect 1928 1102 1933 1103
rect 1938 1102 1943 1103
rect 2952 1103 2954 1107
rect 2954 1103 2957 1107
rect 2962 1103 2965 1107
rect 2965 1103 2967 1107
rect 2952 1102 2957 1103
rect 2962 1102 2967 1103
rect 3976 1103 3978 1107
rect 3978 1103 3981 1107
rect 3986 1103 3989 1107
rect 3989 1103 3991 1107
rect 3976 1102 3981 1103
rect 3986 1102 3991 1103
rect 4285 1087 4290 1092
rect 1437 1067 1442 1072
rect 4173 1037 4178 1042
rect 4269 1027 4274 1032
rect 4189 1007 4194 1012
rect 392 1003 394 1007
rect 394 1003 397 1007
rect 402 1003 405 1007
rect 405 1003 407 1007
rect 392 1002 397 1003
rect 402 1002 407 1003
rect 1416 1003 1418 1007
rect 1418 1003 1421 1007
rect 1426 1003 1429 1007
rect 1429 1003 1431 1007
rect 1416 1002 1421 1003
rect 1426 1002 1431 1003
rect 2440 1003 2442 1007
rect 2442 1003 2445 1007
rect 2450 1003 2453 1007
rect 2453 1003 2455 1007
rect 2440 1002 2445 1003
rect 2450 1002 2455 1003
rect 3472 1003 3474 1007
rect 3474 1003 3477 1007
rect 3482 1003 3485 1007
rect 3485 1003 3487 1007
rect 3472 1002 3477 1003
rect 3482 1002 3487 1003
rect 2541 977 2546 982
rect 1501 967 1506 972
rect 1869 967 1874 972
rect 1501 947 1506 952
rect 1533 907 1538 912
rect 1869 907 1874 912
rect 896 903 898 907
rect 898 903 901 907
rect 906 903 909 907
rect 909 903 911 907
rect 896 902 901 903
rect 906 902 911 903
rect 1928 903 1930 907
rect 1930 903 1933 907
rect 1938 903 1941 907
rect 1941 903 1943 907
rect 1928 902 1933 903
rect 1938 902 1943 903
rect 2952 903 2954 907
rect 2954 903 2957 907
rect 2962 903 2965 907
rect 2965 903 2967 907
rect 2952 902 2957 903
rect 2962 902 2967 903
rect 3976 903 3978 907
rect 3978 903 3981 907
rect 3986 903 3989 907
rect 3989 903 3991 907
rect 3976 902 3981 903
rect 3986 902 3991 903
rect 4141 877 4146 882
rect 392 803 394 807
rect 394 803 397 807
rect 402 803 405 807
rect 405 803 407 807
rect 392 802 397 803
rect 402 802 407 803
rect 1416 803 1418 807
rect 1418 803 1421 807
rect 1426 803 1429 807
rect 1429 803 1431 807
rect 1416 802 1421 803
rect 1426 802 1431 803
rect 2440 803 2442 807
rect 2442 803 2445 807
rect 2450 803 2453 807
rect 2453 803 2455 807
rect 2440 802 2445 803
rect 2450 802 2455 803
rect 3472 803 3474 807
rect 3474 803 3477 807
rect 3482 803 3485 807
rect 3485 803 3487 807
rect 3472 802 3477 803
rect 3482 802 3487 803
rect 1517 797 1522 802
rect 1693 797 1698 802
rect 2061 777 2066 782
rect 2061 757 2066 762
rect 4093 747 4098 752
rect 896 703 898 707
rect 898 703 901 707
rect 906 703 909 707
rect 909 703 911 707
rect 896 702 901 703
rect 906 702 911 703
rect 1928 703 1930 707
rect 1930 703 1933 707
rect 1938 703 1941 707
rect 1941 703 1943 707
rect 1928 702 1933 703
rect 1938 702 1943 703
rect 2952 703 2954 707
rect 2954 703 2957 707
rect 2962 703 2965 707
rect 2965 703 2967 707
rect 2952 702 2957 703
rect 2962 702 2967 703
rect 3976 703 3978 707
rect 3978 703 3981 707
rect 3986 703 3989 707
rect 3989 703 3991 707
rect 3976 702 3981 703
rect 3986 702 3991 703
rect 4077 657 4082 662
rect 392 603 394 607
rect 394 603 397 607
rect 402 603 405 607
rect 405 603 407 607
rect 392 602 397 603
rect 402 602 407 603
rect 1416 603 1418 607
rect 1418 603 1421 607
rect 1426 603 1429 607
rect 1429 603 1431 607
rect 1416 602 1421 603
rect 1426 602 1431 603
rect 2440 603 2442 607
rect 2442 603 2445 607
rect 2450 603 2453 607
rect 2453 603 2455 607
rect 2440 602 2445 603
rect 2450 602 2455 603
rect 3472 603 3474 607
rect 3474 603 3477 607
rect 3482 603 3485 607
rect 3485 603 3487 607
rect 3472 602 3477 603
rect 3482 602 3487 603
rect 896 503 898 507
rect 898 503 901 507
rect 906 503 909 507
rect 909 503 911 507
rect 896 502 901 503
rect 906 502 911 503
rect 1928 503 1930 507
rect 1930 503 1933 507
rect 1938 503 1941 507
rect 1941 503 1943 507
rect 1928 502 1933 503
rect 1938 502 1943 503
rect 2952 503 2954 507
rect 2954 503 2957 507
rect 2962 503 2965 507
rect 2965 503 2967 507
rect 2952 502 2957 503
rect 2962 502 2967 503
rect 3976 503 3978 507
rect 3978 503 3981 507
rect 3986 503 3989 507
rect 3989 503 3991 507
rect 3976 502 3981 503
rect 3986 502 3991 503
rect 4349 477 4354 482
rect 3997 427 4002 432
rect 2541 407 2546 412
rect 392 403 394 407
rect 394 403 397 407
rect 402 403 405 407
rect 405 403 407 407
rect 392 402 397 403
rect 402 402 407 403
rect 1416 403 1418 407
rect 1418 403 1421 407
rect 1426 403 1429 407
rect 1429 403 1431 407
rect 1416 402 1421 403
rect 1426 402 1431 403
rect 2440 403 2442 407
rect 2442 403 2445 407
rect 2450 403 2453 407
rect 2453 403 2455 407
rect 2440 402 2445 403
rect 2450 402 2455 403
rect 3472 403 3474 407
rect 3474 403 3477 407
rect 3482 403 3485 407
rect 3485 403 3487 407
rect 3472 402 3477 403
rect 3482 402 3487 403
rect 3053 397 3058 402
rect 3949 357 3954 362
rect 896 303 898 307
rect 898 303 901 307
rect 906 303 909 307
rect 909 303 911 307
rect 896 302 901 303
rect 906 302 911 303
rect 1928 303 1930 307
rect 1930 303 1933 307
rect 1938 303 1941 307
rect 1941 303 1943 307
rect 1928 302 1933 303
rect 1938 302 1943 303
rect 2952 303 2954 307
rect 2954 303 2957 307
rect 2962 303 2965 307
rect 2965 303 2967 307
rect 2952 302 2957 303
rect 2962 302 2967 303
rect 3976 303 3978 307
rect 3978 303 3981 307
rect 3986 303 3989 307
rect 3989 303 3991 307
rect 3976 302 3981 303
rect 3986 302 3991 303
rect 3949 277 3954 282
rect 4085 267 4090 272
rect 1229 227 1234 232
rect 392 203 394 207
rect 394 203 397 207
rect 402 203 405 207
rect 405 203 407 207
rect 392 202 397 203
rect 402 202 407 203
rect 1416 203 1418 207
rect 1418 203 1421 207
rect 1426 203 1429 207
rect 1429 203 1431 207
rect 1416 202 1421 203
rect 1426 202 1431 203
rect 2440 203 2442 207
rect 2442 203 2445 207
rect 2450 203 2453 207
rect 2453 203 2455 207
rect 2440 202 2445 203
rect 2450 202 2455 203
rect 3472 203 3474 207
rect 3474 203 3477 207
rect 3482 203 3485 207
rect 3485 203 3487 207
rect 3472 202 3477 203
rect 3482 202 3487 203
rect 4237 157 4242 162
rect 4381 157 4386 162
rect 4365 147 4370 152
rect 4301 127 4306 132
rect 4317 127 4322 132
rect 4221 107 4226 112
rect 896 103 898 107
rect 898 103 901 107
rect 906 103 909 107
rect 909 103 911 107
rect 896 102 901 103
rect 906 102 911 103
rect 1928 103 1930 107
rect 1930 103 1933 107
rect 1938 103 1941 107
rect 1941 103 1943 107
rect 1928 102 1933 103
rect 1938 102 1943 103
rect 2952 103 2954 107
rect 2954 103 2957 107
rect 2962 103 2965 107
rect 2965 103 2967 107
rect 2952 102 2957 103
rect 2962 102 2967 103
rect 3976 103 3978 107
rect 3978 103 3981 107
rect 3986 103 3989 107
rect 3989 103 3991 107
rect 3976 102 3981 103
rect 3986 102 3991 103
rect 4125 97 4130 102
rect 4141 87 4146 92
rect 4205 87 4210 92
rect 4333 67 4338 72
rect 4157 37 4162 42
rect 392 3 394 7
rect 394 3 397 7
rect 402 3 405 7
rect 405 3 407 7
rect 392 2 397 3
rect 402 2 407 3
rect 1416 3 1418 7
rect 1418 3 1421 7
rect 1426 3 1429 7
rect 1429 3 1431 7
rect 1416 2 1421 3
rect 1426 2 1431 3
rect 2440 3 2442 7
rect 2442 3 2445 7
rect 2450 3 2453 7
rect 2453 3 2455 7
rect 2440 2 2445 3
rect 2450 2 2455 3
rect 3472 3 3474 7
rect 3474 3 3477 7
rect 3482 3 3485 7
rect 3485 3 3487 7
rect 3472 2 3477 3
rect 3482 2 3487 3
<< metal6 >>
rect 392 3007 408 3130
rect 397 3002 402 3007
rect 407 3002 408 3007
rect 392 2807 408 3002
rect 397 2802 402 2807
rect 407 2802 408 2807
rect 392 2607 408 2802
rect 397 2602 402 2607
rect 407 2602 408 2607
rect 392 2407 408 2602
rect 397 2402 402 2407
rect 407 2402 408 2407
rect 392 2207 408 2402
rect 397 2202 402 2207
rect 407 2202 408 2207
rect 392 2007 408 2202
rect 397 2002 402 2007
rect 407 2002 408 2007
rect 392 1807 408 2002
rect 397 1802 402 1807
rect 407 1802 408 1807
rect 392 1607 408 1802
rect 397 1602 402 1607
rect 407 1602 408 1607
rect 392 1407 408 1602
rect 397 1402 402 1407
rect 407 1402 408 1407
rect 392 1207 408 1402
rect 397 1202 402 1207
rect 407 1202 408 1207
rect 392 1007 408 1202
rect 397 1002 402 1007
rect 407 1002 408 1007
rect 392 807 408 1002
rect 397 802 402 807
rect 407 802 408 807
rect 392 607 408 802
rect 397 602 402 607
rect 407 602 408 607
rect 392 407 408 602
rect 397 402 402 407
rect 407 402 408 407
rect 392 207 408 402
rect 397 202 402 207
rect 407 202 408 207
rect 392 7 408 202
rect 397 2 402 7
rect 407 2 408 7
rect 392 -30 408 2
rect 896 3107 912 3130
rect 901 3102 906 3107
rect 911 3102 912 3107
rect 896 2907 912 3102
rect 901 2902 906 2907
rect 911 2902 912 2907
rect 896 2707 912 2902
rect 901 2702 906 2707
rect 911 2702 912 2707
rect 896 2507 912 2702
rect 901 2502 906 2507
rect 911 2502 912 2507
rect 896 2307 912 2502
rect 901 2302 906 2307
rect 911 2302 912 2307
rect 896 2107 912 2302
rect 901 2102 906 2107
rect 911 2102 912 2107
rect 896 1907 912 2102
rect 901 1902 906 1907
rect 911 1902 912 1907
rect 896 1707 912 1902
rect 901 1702 906 1707
rect 911 1702 912 1707
rect 896 1507 912 1702
rect 901 1502 906 1507
rect 911 1502 912 1507
rect 896 1307 912 1502
rect 901 1302 906 1307
rect 911 1302 912 1307
rect 896 1107 912 1302
rect 1416 3007 1432 3130
rect 1421 3002 1426 3007
rect 1431 3002 1432 3007
rect 1416 2807 1432 3002
rect 1421 2802 1426 2807
rect 1431 2802 1432 2807
rect 1416 2607 1432 2802
rect 1421 2602 1426 2607
rect 1431 2602 1432 2607
rect 1416 2407 1432 2602
rect 1421 2402 1426 2407
rect 1431 2402 1432 2407
rect 1416 2207 1432 2402
rect 1928 3107 1944 3130
rect 1933 3102 1938 3107
rect 1943 3102 1944 3107
rect 1928 2907 1944 3102
rect 1933 2902 1938 2907
rect 1943 2902 1944 2907
rect 1928 2707 1944 2902
rect 1933 2702 1938 2707
rect 1943 2702 1944 2707
rect 1928 2507 1944 2702
rect 1933 2502 1938 2507
rect 1943 2502 1944 2507
rect 1869 2322 1874 2347
rect 1421 2202 1426 2207
rect 1431 2202 1432 2207
rect 1416 2007 1432 2202
rect 1928 2307 1944 2502
rect 2440 3007 2456 3130
rect 2445 3002 2450 3007
rect 2455 3002 2456 3007
rect 2440 2807 2456 3002
rect 2445 2802 2450 2807
rect 2455 2802 2456 2807
rect 2440 2607 2456 2802
rect 2445 2602 2450 2607
rect 2455 2602 2456 2607
rect 1933 2302 1938 2307
rect 1943 2302 1944 2307
rect 1928 2107 1944 2302
rect 1933 2102 1938 2107
rect 1943 2102 1944 2107
rect 1421 2002 1426 2007
rect 1431 2002 1432 2007
rect 1416 1807 1432 2002
rect 1421 1802 1426 1807
rect 1431 1802 1432 1807
rect 1416 1607 1432 1802
rect 1421 1602 1426 1607
rect 1431 1602 1432 1607
rect 1416 1407 1432 1602
rect 1421 1402 1426 1407
rect 1431 1402 1432 1407
rect 1416 1207 1432 1402
rect 1421 1202 1426 1207
rect 1431 1202 1432 1207
rect 901 1102 906 1107
rect 911 1102 912 1107
rect 896 907 912 1102
rect 901 902 906 907
rect 911 902 912 907
rect 896 707 912 902
rect 901 702 906 707
rect 911 702 912 707
rect 896 507 912 702
rect 901 502 906 507
rect 911 502 912 507
rect 896 307 912 502
rect 901 302 906 307
rect 911 302 912 307
rect 896 107 912 302
rect 1229 232 1234 1127
rect 1416 1007 1432 1202
rect 1437 1072 1442 1597
rect 1421 1002 1426 1007
rect 1431 1002 1432 1007
rect 1416 807 1432 1002
rect 1501 952 1506 967
rect 1421 802 1426 807
rect 1431 802 1432 807
rect 1416 607 1432 802
rect 1517 802 1522 1337
rect 1533 1202 1538 1247
rect 1549 1232 1554 1317
rect 1581 1132 1586 1447
rect 1613 1182 1618 1857
rect 1533 912 1538 1127
rect 1693 802 1698 1467
rect 1725 1182 1730 2067
rect 1789 1312 1794 1327
rect 1837 1302 1842 1317
rect 1901 1222 1906 1937
rect 1928 1907 1944 2102
rect 1933 1902 1938 1907
rect 1943 1902 1944 1907
rect 1928 1707 1944 1902
rect 1933 1702 1938 1707
rect 1943 1702 1944 1707
rect 1928 1507 1944 1702
rect 1997 2352 2002 2427
rect 1997 1592 2002 2347
rect 2440 2407 2456 2602
rect 2952 3107 2968 3130
rect 2957 3102 2962 3107
rect 2967 3102 2968 3107
rect 2952 2907 2968 3102
rect 2957 2902 2962 2907
rect 2967 2902 2968 2907
rect 2952 2707 2968 2902
rect 3472 3007 3488 3130
rect 3477 3002 3482 3007
rect 3487 3002 3488 3007
rect 3472 2807 3488 3002
rect 3477 2802 3482 2807
rect 3487 2802 3488 2807
rect 2957 2702 2962 2707
rect 2967 2702 2968 2707
rect 2952 2507 2968 2702
rect 2957 2502 2962 2507
rect 2967 2502 2968 2507
rect 2941 2472 2946 2497
rect 2445 2402 2450 2407
rect 2455 2402 2456 2407
rect 2440 2207 2456 2402
rect 2445 2202 2450 2207
rect 2455 2202 2456 2207
rect 2440 2007 2456 2202
rect 2445 2002 2450 2007
rect 2455 2002 2456 2007
rect 2440 1807 2456 2002
rect 2445 1802 2450 1807
rect 2455 1802 2456 1807
rect 2205 1712 2210 1747
rect 2440 1607 2456 1802
rect 2445 1602 2450 1607
rect 2455 1602 2456 1607
rect 1933 1502 1938 1507
rect 1943 1502 1944 1507
rect 1928 1307 1944 1502
rect 2429 1412 2434 1427
rect 2440 1407 2456 1602
rect 1933 1302 1938 1307
rect 1943 1302 1944 1307
rect 1928 1107 1944 1302
rect 2445 1402 2450 1407
rect 2455 1402 2456 1407
rect 2440 1207 2456 1402
rect 2952 2307 2968 2502
rect 2957 2302 2962 2307
rect 2967 2302 2968 2307
rect 2952 2107 2968 2302
rect 2957 2102 2962 2107
rect 2967 2102 2968 2107
rect 2952 1907 2968 2102
rect 2957 1902 2962 1907
rect 2967 1902 2968 1907
rect 2952 1707 2968 1902
rect 2957 1702 2962 1707
rect 2967 1702 2968 1707
rect 2952 1507 2968 1702
rect 2957 1502 2962 1507
rect 2967 1502 2968 1507
rect 2952 1307 2968 1502
rect 2957 1302 2962 1307
rect 2967 1302 2968 1307
rect 2941 1252 2946 1277
rect 2445 1202 2450 1207
rect 2455 1202 2456 1207
rect 2189 1142 2194 1157
rect 1933 1102 1938 1107
rect 1943 1102 1944 1107
rect 1869 912 1874 967
rect 1928 907 1944 1102
rect 1933 902 1938 907
rect 1943 902 1944 907
rect 1421 602 1426 607
rect 1431 602 1432 607
rect 1416 407 1432 602
rect 1421 402 1426 407
rect 1431 402 1432 407
rect 901 102 906 107
rect 911 102 912 107
rect 896 -30 912 102
rect 1416 207 1432 402
rect 1421 202 1426 207
rect 1431 202 1432 207
rect 1416 7 1432 202
rect 1421 2 1426 7
rect 1431 2 1432 7
rect 1416 -30 1432 2
rect 1928 707 1944 902
rect 2440 1007 2456 1202
rect 2445 1002 2450 1007
rect 2455 1002 2456 1007
rect 2440 807 2456 1002
rect 2952 1107 2968 1302
rect 3101 1152 3106 2467
rect 3197 1212 3202 2757
rect 3472 2607 3488 2802
rect 3477 2602 3482 2607
rect 3487 2602 3488 2607
rect 3472 2407 3488 2602
rect 3477 2402 3482 2407
rect 3487 2402 3488 2407
rect 3472 2207 3488 2402
rect 3477 2202 3482 2207
rect 3487 2202 3488 2207
rect 3277 2052 3282 2187
rect 3472 2007 3488 2202
rect 3477 2002 3482 2007
rect 3487 2002 3488 2007
rect 3472 1807 3488 2002
rect 3477 1802 3482 1807
rect 3487 1802 3488 1807
rect 3472 1607 3488 1802
rect 3477 1602 3482 1607
rect 3487 1602 3488 1607
rect 3472 1407 3488 1602
rect 3477 1402 3482 1407
rect 3487 1402 3488 1407
rect 3472 1207 3488 1402
rect 3477 1202 3482 1207
rect 3487 1202 3488 1207
rect 2957 1102 2962 1107
rect 2967 1102 2968 1107
rect 2445 802 2450 807
rect 2455 802 2456 807
rect 2061 762 2066 777
rect 1933 702 1938 707
rect 1943 702 1944 707
rect 1928 507 1944 702
rect 1933 502 1938 507
rect 1943 502 1944 507
rect 1928 307 1944 502
rect 1933 302 1938 307
rect 1943 302 1944 307
rect 1928 107 1944 302
rect 1933 102 1938 107
rect 1943 102 1944 107
rect 1928 -30 1944 102
rect 2440 607 2456 802
rect 2445 602 2450 607
rect 2455 602 2456 607
rect 2440 407 2456 602
rect 2541 412 2546 977
rect 2952 907 2968 1102
rect 2957 902 2962 907
rect 2967 902 2968 907
rect 2952 707 2968 902
rect 2957 702 2962 707
rect 2967 702 2968 707
rect 2952 507 2968 702
rect 2957 502 2962 507
rect 2967 502 2968 507
rect 2445 402 2450 407
rect 2455 402 2456 407
rect 2440 207 2456 402
rect 2445 202 2450 207
rect 2455 202 2456 207
rect 2440 7 2456 202
rect 2445 2 2450 7
rect 2455 2 2456 7
rect 2440 -30 2456 2
rect 2952 307 2968 502
rect 3053 402 3058 1127
rect 3472 1007 3488 1202
rect 3477 1002 3482 1007
rect 3487 1002 3488 1007
rect 3472 807 3488 1002
rect 3477 802 3482 807
rect 3487 802 3488 807
rect 3472 607 3488 802
rect 3477 602 3482 607
rect 3487 602 3488 607
rect 3472 407 3488 602
rect 3477 402 3482 407
rect 3487 402 3488 407
rect 2957 302 2962 307
rect 2967 302 2968 307
rect 2952 107 2968 302
rect 2957 102 2962 107
rect 2967 102 2968 107
rect 2952 -30 2968 102
rect 3472 207 3488 402
rect 3976 3107 3992 3130
rect 3981 3102 3986 3107
rect 3991 3102 3992 3107
rect 3976 2907 3992 3102
rect 3981 2902 3986 2907
rect 3991 2902 3992 2907
rect 3976 2707 3992 2902
rect 3981 2702 3986 2707
rect 3991 2702 3992 2707
rect 3976 2507 3992 2702
rect 3981 2502 3986 2507
rect 3991 2502 3992 2507
rect 3976 2307 3992 2502
rect 3981 2302 3986 2307
rect 3991 2302 3992 2307
rect 3976 2107 3992 2302
rect 3981 2102 3986 2107
rect 3991 2102 3992 2107
rect 3976 1907 3992 2102
rect 3981 1902 3986 1907
rect 3991 1902 3992 1907
rect 3976 1707 3992 1902
rect 3981 1702 3986 1707
rect 3991 1702 3992 1707
rect 3976 1507 3992 1702
rect 3981 1502 3986 1507
rect 3991 1502 3992 1507
rect 3976 1307 3992 1502
rect 3981 1302 3986 1307
rect 3991 1302 3992 1307
rect 3976 1107 3992 1302
rect 3981 1102 3986 1107
rect 3991 1102 3992 1107
rect 3976 907 3992 1102
rect 3981 902 3986 907
rect 3991 902 3992 907
rect 3976 707 3992 902
rect 3981 702 3986 707
rect 3991 702 3992 707
rect 3976 507 3992 702
rect 3981 502 3986 507
rect 3991 502 3992 507
rect 3949 282 3954 357
rect 3976 307 3992 502
rect 3997 432 4002 1847
rect 4077 1272 4082 2147
rect 4093 752 4098 2147
rect 3981 302 3986 307
rect 3991 302 3992 307
rect 3477 202 3482 207
rect 3487 202 3488 207
rect 3472 7 3488 202
rect 3477 2 3482 7
rect 3487 2 3488 7
rect 3472 -30 3488 2
rect 3976 107 3992 302
rect 4077 272 4082 657
rect 4077 267 4085 272
rect 3981 102 3986 107
rect 3991 102 3992 107
rect 3976 -30 3992 102
rect 4125 102 4130 2767
rect 4141 92 4146 877
rect 4157 42 4162 1567
rect 4173 1042 4178 1727
rect 4189 1012 4194 1937
rect 4205 92 4210 1697
rect 4221 112 4226 1277
rect 4237 162 4242 2017
rect 4253 1782 4258 3047
rect 4269 1032 4274 3037
rect 4301 2652 4306 3067
rect 4285 1092 4290 1787
rect 4301 1122 4306 2347
rect 4301 132 4306 1107
rect 4317 132 4322 2737
rect 4333 72 4338 1817
rect 4349 1802 4354 2747
rect 4349 482 4354 1787
rect 4365 152 4370 2437
rect 4381 162 4386 2357
use BUFX2  BUFX2_40
timestamp 1751266522
transform -1 0 28 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_52
timestamp 1751266522
transform -1 0 52 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_81
timestamp 1751266522
transform -1 0 228 0 -1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_57
timestamp 1751266522
transform 1 0 4 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_50
timestamp 1751266522
transform 1 0 76 0 1 105
box -2 -3 74 103
use DFFSR  DFFSR_21
timestamp 1751266522
transform 1 0 148 0 1 105
box -2 -3 178 103
use BUFX2  BUFX2_60
timestamp 1751266522
transform 1 0 228 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_66
timestamp 1751266522
transform 1 0 252 0 -1 105
box -2 -3 74 103
use BUFX2  BUFX2_24
timestamp 1751266522
transform -1 0 348 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_22
timestamp 1751266522
transform 1 0 348 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_29
timestamp 1751266522
transform -1 0 348 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_56
timestamp 1751266522
transform -1 0 372 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_54
timestamp 1751266522
transform 1 0 372 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1751266522
transform 1 0 396 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1751266522
transform 1 0 404 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_59
timestamp 1751266522
transform 1 0 412 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_83
timestamp 1751266522
transform -1 0 612 0 -1 105
box -2 -3 178 103
use FILL  FILL_1_0_0
timestamp 1751266522
transform -1 0 380 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1751266522
transform -1 0 388 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_85
timestamp 1751266522
transform -1 0 564 0 1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_149
timestamp 1751266522
transform -1 0 644 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_26
timestamp 1751266522
transform 1 0 644 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_17
timestamp 1751266522
transform 1 0 668 0 -1 105
box -2 -3 178 103
use BUFX2  BUFX2_53
timestamp 1751266522
transform -1 0 588 0 1 105
box -2 -3 26 103
use DFFSR  DFFSR_82
timestamp 1751266522
transform -1 0 764 0 1 105
box -2 -3 178 103
use BUFX2  BUFX2_23
timestamp 1751266522
transform -1 0 788 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_146
timestamp 1751266522
transform -1 0 820 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_18
timestamp 1751266522
transform 1 0 820 0 1 105
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1751266522
transform -1 0 884 0 1 105
box -2 -3 18 103
use INVX1  INVX1_9
timestamp 1751266522
transform 1 0 852 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_148
timestamp 1751266522
transform -1 0 876 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1751266522
transform 1 0 884 0 1 105
box -2 -3 34 103
use FILL  FILL_0_1_1
timestamp 1751266522
transform 1 0 908 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_0
timestamp 1751266522
transform 1 0 900 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_25
timestamp 1751266522
transform 1 0 876 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_11
timestamp 1751266522
transform 1 0 932 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_1
timestamp 1751266522
transform 1 0 924 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_0
timestamp 1751266522
transform 1 0 916 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_142
timestamp 1751266522
transform 1 0 916 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1751266522
transform 1 0 964 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_21
timestamp 1751266522
transform 1 0 972 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_19
timestamp 1751266522
transform 1 0 948 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_31
timestamp 1751266522
transform 1 0 996 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_144
timestamp 1751266522
transform 1 0 996 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1751266522
transform 1 0 1028 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_143
timestamp 1751266522
transform 1 0 1028 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1751266522
transform 1 0 1076 0 1 105
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1751266522
transform 1 0 1060 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_16
timestamp 1751266522
transform -1 0 1108 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_20
timestamp 1751266522
transform 1 0 1060 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_9
timestamp 1751266522
transform -1 0 1132 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_10
timestamp 1751266522
transform -1 0 1148 0 -1 105
box -2 -3 18 103
use DFFSR  DFFSR_19
timestamp 1751266522
transform 1 0 1148 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_20
timestamp 1751266522
transform 1 0 1108 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1751266522
transform 1 0 1140 0 1 105
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1751266522
transform 1 0 1172 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_22
timestamp 1751266522
transform 1 0 1188 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1751266522
transform 1 0 1220 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1751266522
transform 1 0 1252 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1751266522
transform 1 0 1348 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_25
timestamp 1751266522
transform 1 0 1316 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1751266522
transform 1 0 1284 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_57
timestamp 1751266522
transform -1 0 1372 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1751266522
transform 1 0 1324 0 -1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_6
timestamp 1751266522
transform 1 0 1436 0 1 105
box -2 -3 42 103
use FILL  FILL_1_2_1
timestamp 1751266522
transform 1 0 1428 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_0
timestamp 1751266522
transform 1 0 1420 0 1 105
box -2 -3 10 103
use NAND3X1  NAND3X1_72
timestamp 1751266522
transform -1 0 1420 0 1 105
box -2 -3 34 103
use FILL  FILL_0_2_1
timestamp 1751266522
transform 1 0 1428 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_0
timestamp 1751266522
transform 1 0 1420 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_10
timestamp 1751266522
transform 1 0 1396 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_13
timestamp 1751266522
transform 1 0 1372 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_203
timestamp 1751266522
transform 1 0 1436 0 -1 105
box -2 -3 178 103
use DFFSR  DFFSR_165
timestamp 1751266522
transform -1 0 1788 0 -1 105
box -2 -3 178 103
use NAND3X1  NAND3X1_74
timestamp 1751266522
transform -1 0 1508 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_53
timestamp 1751266522
transform -1 0 1532 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_51
timestamp 1751266522
transform -1 0 1556 0 1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_5
timestamp 1751266522
transform 1 0 1556 0 1 105
box -2 -3 42 103
use AOI22X1  AOI22X1_1
timestamp 1751266522
transform 1 0 1596 0 1 105
box -2 -3 42 103
use DFFSR  DFFSR_133
timestamp 1751266522
transform -1 0 1964 0 -1 105
box -2 -3 178 103
use DFFSR  DFFSR_134
timestamp 1751266522
transform -1 0 1812 0 1 105
box -2 -3 178 103
use INVX2  INVX2_93
timestamp 1751266522
transform 1 0 1812 0 1 105
box -2 -3 18 103
use INVX8  INVX8_21
timestamp 1751266522
transform -1 0 1868 0 1 105
box -2 -3 42 103
use OAI22X1  OAI22X1_111
timestamp 1751266522
transform 1 0 1900 0 1 105
box -2 -3 42 103
use BUFX4  BUFX4_165
timestamp 1751266522
transform 1 0 1868 0 1 105
box -2 -3 34 103
use FILL  FILL_1_3_1
timestamp 1751266522
transform -1 0 1956 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_0
timestamp 1751266522
transform -1 0 1948 0 1 105
box -2 -3 10 103
use INVX1  INVX1_156
timestamp 1751266522
transform -1 0 2004 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_622
timestamp 1751266522
transform -1 0 1988 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1751266522
transform 1 0 1980 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_3_1
timestamp 1751266522
transform 1 0 1972 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_0
timestamp 1751266522
transform 1 0 1964 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_542
timestamp 1751266522
transform 1 0 2052 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_179
timestamp 1751266522
transform 1 0 2020 0 1 105
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1751266522
transform 1 0 2004 0 1 105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_24
timestamp 1751266522
transform 1 0 2060 0 -1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_176
timestamp 1751266522
transform -1 0 2060 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_227
timestamp 1751266522
transform 1 0 2012 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_231
timestamp 1751266522
transform 1 0 2148 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_543
timestamp 1751266522
transform 1 0 2116 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_544
timestamp 1751266522
transform -1 0 2116 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_174
timestamp 1751266522
transform -1 0 2156 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_621
timestamp 1751266522
transform -1 0 2204 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_170
timestamp 1751266522
transform 1 0 2156 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_189
timestamp 1751266522
transform -1 0 2212 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_187
timestamp 1751266522
transform 1 0 2212 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_190
timestamp 1751266522
transform -1 0 2276 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_185
timestamp 1751266522
transform -1 0 2308 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1751266522
transform -1 0 2332 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_188
timestamp 1751266522
transform 1 0 2332 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_186
timestamp 1751266522
transform 1 0 2204 0 1 105
box -2 -3 34 103
use INVX2  INVX2_146
timestamp 1751266522
transform -1 0 2252 0 1 105
box -2 -3 18 103
use DFFSR  DFFSR_164
timestamp 1751266522
transform -1 0 2428 0 1 105
box -2 -3 178 103
use FILL  FILL_1_4_0
timestamp 1751266522
transform 1 0 2444 0 1 105
box -2 -3 10 103
use INVX2  INVX2_122
timestamp 1751266522
transform 1 0 2428 0 1 105
box -2 -3 18 103
use FILL  FILL_0_4_1
timestamp 1751266522
transform -1 0 2436 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_4_0
timestamp 1751266522
transform -1 0 2428 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_247
timestamp 1751266522
transform -1 0 2420 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_184
timestamp 1751266522
transform 1 0 2364 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_546
timestamp 1751266522
transform -1 0 2564 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_181
timestamp 1751266522
transform -1 0 2532 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_73
timestamp 1751266522
transform 1 0 2460 0 1 105
box -2 -3 42 103
use FILL  FILL_1_4_1
timestamp 1751266522
transform 1 0 2452 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_166
timestamp 1751266522
transform -1 0 2612 0 -1 105
box -2 -3 178 103
use AOI21X1  AOI21X1_174
timestamp 1751266522
transform -1 0 2644 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_534
timestamp 1751266522
transform -1 0 2676 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_535
timestamp 1751266522
transform 1 0 2676 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_175
timestamp 1751266522
transform 1 0 2708 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_177
timestamp 1751266522
transform 1 0 2564 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_539
timestamp 1751266522
transform -1 0 2628 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_72
timestamp 1751266522
transform -1 0 2668 0 1 105
box -2 -3 42 103
use AOI21X1  AOI21X1_178
timestamp 1751266522
transform -1 0 2700 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1751266522
transform -1 0 2732 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_71
timestamp 1751266522
transform -1 0 2780 0 -1 105
box -2 -3 42 103
use DFFSR  DFFSR_168
timestamp 1751266522
transform -1 0 2956 0 -1 105
box -2 -3 178 103
use NAND2X1  NAND2X1_256
timestamp 1751266522
transform 1 0 2732 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_700
timestamp 1751266522
transform -1 0 2788 0 1 105
box -2 -3 34 103
use DFFSR  DFFSR_139
timestamp 1751266522
transform 1 0 2788 0 1 105
box -2 -3 178 103
use FILL  FILL_0_5_0
timestamp 1751266522
transform 1 0 2956 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1751266522
transform 1 0 2964 0 -1 105
box -2 -3 10 103
use INVX2  INVX2_91
timestamp 1751266522
transform 1 0 2972 0 -1 105
box -2 -3 18 103
use DFFSR  DFFSR_197
timestamp 1751266522
transform -1 0 3164 0 -1 105
box -2 -3 178 103
use FILL  FILL_1_5_0
timestamp 1751266522
transform -1 0 2972 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_1
timestamp 1751266522
transform -1 0 2980 0 1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_52
timestamp 1751266522
transform -1 0 3052 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_20
timestamp 1751266522
transform 1 0 3052 0 1 105
box -2 -3 74 103
use OAI21X1  OAI21X1_459
timestamp 1751266522
transform 1 0 3164 0 -1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_65
timestamp 1751266522
transform 1 0 3196 0 -1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_460
timestamp 1751266522
transform 1 0 3236 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_45
timestamp 1751266522
transform -1 0 3196 0 1 105
box -2 -3 74 103
use DFFSR  DFFSR_210
timestamp 1751266522
transform -1 0 3372 0 1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_63
timestamp 1751266522
transform -1 0 3340 0 -1 105
box -2 -3 74 103
use DFFSR  DFFSR_228
timestamp 1751266522
transform -1 0 3516 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_458
timestamp 1751266522
transform -1 0 3404 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_148
timestamp 1751266522
transform 1 0 3404 0 1 105
box -2 -3 34 103
use FILL  FILL_1_6_0
timestamp 1751266522
transform -1 0 3444 0 1 105
box -2 -3 10 103
use FILL  FILL_0_6_0
timestamp 1751266522
transform 1 0 3516 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_6_1
timestamp 1751266522
transform 1 0 3524 0 -1 105
box -2 -3 10 103
use INVX2  INVX2_145
timestamp 1751266522
transform 1 0 3532 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_378
timestamp 1751266522
transform 1 0 3548 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_107
timestamp 1751266522
transform 1 0 3580 0 -1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_48
timestamp 1751266522
transform 1 0 3612 0 -1 105
box -2 -3 42 103
use FILL  FILL_1_6_1
timestamp 1751266522
transform -1 0 3452 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_196
timestamp 1751266522
transform -1 0 3628 0 1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_376
timestamp 1751266522
transform -1 0 3684 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_105
timestamp 1751266522
transform 1 0 3684 0 -1 105
box -2 -3 34 103
use DFFSR  DFFSR_198
timestamp 1751266522
transform -1 0 3892 0 -1 105
box -2 -3 178 103
use DFFSR  DFFSR_230
timestamp 1751266522
transform -1 0 3804 0 1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_377
timestamp 1751266522
transform 1 0 3804 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_104
timestamp 1751266522
transform -1 0 3900 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_106
timestamp 1751266522
transform 1 0 3836 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_47
timestamp 1751266522
transform -1 0 3972 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_375
timestamp 1751266522
transform -1 0 3932 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_10
timestamp 1751266522
transform -1 0 3964 0 -1 105
box -2 -3 74 103
use FILL  FILL_1_7_1
timestamp 1751266522
transform 1 0 3980 0 1 105
box -2 -3 10 103
use FILL  FILL_1_7_0
timestamp 1751266522
transform 1 0 3972 0 1 105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_53
timestamp 1751266522
transform 1 0 3980 0 -1 105
box -2 -3 74 103
use FILL  FILL_0_7_1
timestamp 1751266522
transform 1 0 3972 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_7_0
timestamp 1751266522
transform 1 0 3964 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_68
timestamp 1751266522
transform 1 0 4052 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_138
timestamp 1751266522
transform -1 0 4108 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_83
timestamp 1751266522
transform -1 0 4140 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_206
timestamp 1751266522
transform 1 0 4140 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_123
timestamp 1751266522
transform 1 0 3988 0 1 105
box -2 -3 18 103
use INVX2  INVX2_92
timestamp 1751266522
transform -1 0 4020 0 1 105
box -2 -3 18 103
use DFFSR  DFFSR_229
timestamp 1751266522
transform -1 0 4196 0 1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_7
timestamp 1751266522
transform -1 0 4268 0 1 105
box -2 -3 74 103
use INVX8  INVX8_13
timestamp 1751266522
transform 1 0 4204 0 -1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_212
timestamp 1751266522
transform -1 0 4204 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1751266522
transform 1 0 4300 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_228
timestamp 1751266522
transform -1 0 4300 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_91
timestamp 1751266522
transform 1 0 4308 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_204
timestamp 1751266522
transform 1 0 4276 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_139
timestamp 1751266522
transform 1 0 4244 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_81
timestamp 1751266522
transform -1 0 4356 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_50
timestamp 1751266522
transform 1 0 4340 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1751266522
transform -1 0 4380 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1751266522
transform -1 0 4388 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_3
timestamp 1751266522
transform -1 0 4396 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_93
timestamp 1751266522
transform -1 0 4380 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1751266522
transform 1 0 4380 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1751266522
transform 1 0 4388 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_69
timestamp 1751266522
transform -1 0 180 0 -1 305
box -2 -3 178 103
use DFFSR  DFFSR_24
timestamp 1751266522
transform 1 0 180 0 -1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_147
timestamp 1751266522
transform -1 0 388 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1751266522
transform 1 0 388 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1751266522
transform 1 0 396 0 -1 305
box -2 -3 10 103
use BUFX2  BUFX2_14
timestamp 1751266522
transform 1 0 404 0 -1 305
box -2 -3 26 103
use DFFSR  DFFSR_88
timestamp 1751266522
transform -1 0 604 0 -1 305
box -2 -3 178 103
use DFFSR  DFFSR_23
timestamp 1751266522
transform 1 0 604 0 -1 305
box -2 -3 178 103
use BUFX2  BUFX2_66
timestamp 1751266522
transform 1 0 780 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_30
timestamp 1751266522
transform 1 0 804 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1751266522
transform 1 0 836 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_32
timestamp 1751266522
transform 1 0 852 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1751266522
transform 1 0 884 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1751266522
transform 1 0 916 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1751266522
transform 1 0 924 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_29
timestamp 1751266522
transform 1 0 932 0 -1 305
box -2 -3 34 103
use DFFSR  DFFSR_18
timestamp 1751266522
transform 1 0 964 0 -1 305
box -2 -3 178 103
use INVX1  INVX1_14
timestamp 1751266522
transform -1 0 1156 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_27
timestamp 1751266522
transform 1 0 1156 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_15
timestamp 1751266522
transform -1 0 1212 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_14
timestamp 1751266522
transform -1 0 1236 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_12
timestamp 1751266522
transform 1 0 1236 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_4
timestamp 1751266522
transform 1 0 1260 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_73
timestamp 1751266522
transform -1 0 1332 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_52
timestamp 1751266522
transform 1 0 1332 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_10
timestamp 1751266522
transform 1 0 1356 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_76
timestamp 1751266522
transform -1 0 1428 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_2_0
timestamp 1751266522
transform 1 0 1428 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1751266522
transform 1 0 1436 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_163
timestamp 1751266522
transform 1 0 1444 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_55
timestamp 1751266522
transform -1 0 1492 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_3
timestamp 1751266522
transform 1 0 1492 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_58
timestamp 1751266522
transform -1 0 1556 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_9
timestamp 1751266522
transform 1 0 1556 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_165
timestamp 1751266522
transform -1 0 1620 0 -1 305
box -2 -3 26 103
use DFFSR  DFFSR_167
timestamp 1751266522
transform -1 0 1796 0 -1 305
box -2 -3 178 103
use AOI22X1  AOI22X1_13
timestamp 1751266522
transform 1 0 1796 0 -1 305
box -2 -3 42 103
use DFFSR  DFFSR_132
timestamp 1751266522
transform -1 0 2012 0 -1 305
box -2 -3 178 103
use FILL  FILL_2_3_0
timestamp 1751266522
transform 1 0 2012 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1751266522
transform 1 0 2020 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_627
timestamp 1751266522
transform 1 0 2028 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_233
timestamp 1751266522
transform 1 0 2060 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_122
timestamp 1751266522
transform 1 0 2084 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_624
timestamp 1751266522
transform -1 0 2132 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_619
timestamp 1751266522
transform -1 0 2164 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_620
timestamp 1751266522
transform 1 0 2164 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1751266522
transform 1 0 2196 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_617
timestamp 1751266522
transform -1 0 2252 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1751266522
transform -1 0 2284 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1751266522
transform -1 0 2308 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_227
timestamp 1751266522
transform 1 0 2308 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_609
timestamp 1751266522
transform -1 0 2364 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_119
timestamp 1751266522
transform 1 0 2364 0 -1 305
box -2 -3 18 103
use BUFX4  BUFX4_1
timestamp 1751266522
transform 1 0 2380 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_528
timestamp 1751266522
transform -1 0 2444 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_4_0
timestamp 1751266522
transform -1 0 2452 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1751266522
transform -1 0 2460 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_529
timestamp 1751266522
transform -1 0 2492 0 -1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_108
timestamp 1751266522
transform 1 0 2492 0 -1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_545
timestamp 1751266522
transform 1 0 2532 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_180
timestamp 1751266522
transform -1 0 2596 0 -1 305
box -2 -3 34 103
use DFFSR  DFFSR_170
timestamp 1751266522
transform -1 0 2772 0 -1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_699
timestamp 1751266522
transform -1 0 2804 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_137
timestamp 1751266522
transform 1 0 2804 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_697
timestamp 1751266522
transform -1 0 2852 0 -1 305
box -2 -3 34 103
use DFFSR  DFFSR_202
timestamp 1751266522
transform -1 0 3028 0 -1 305
box -2 -3 178 103
use FILL  FILL_2_5_0
timestamp 1751266522
transform -1 0 3036 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1751266522
transform -1 0 3044 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_678
timestamp 1751266522
transform -1 0 3076 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_679
timestamp 1751266522
transform 1 0 3076 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_85
timestamp 1751266522
transform 1 0 3108 0 -1 305
box -2 -3 42 103
use DFFSR  DFFSR_232
timestamp 1751266522
transform -1 0 3324 0 -1 305
box -2 -3 178 103
use INVX2  INVX2_136
timestamp 1751266522
transform 1 0 3324 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_369
timestamp 1751266522
transform 1 0 3340 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_145
timestamp 1751266522
transform -1 0 3404 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_244
timestamp 1751266522
transform -1 0 3436 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_249
timestamp 1751266522
transform 1 0 3436 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_6_0
timestamp 1751266522
transform 1 0 3468 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1751266522
transform 1 0 3476 0 -1 305
box -2 -3 10 103
use AOI22X1  AOI22X1_45
timestamp 1751266522
transform 1 0 3484 0 -1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_99
timestamp 1751266522
transform -1 0 3556 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_368
timestamp 1751266522
transform 1 0 3556 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_98
timestamp 1751266522
transform 1 0 3588 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_147
timestamp 1751266522
transform 1 0 3620 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_463
timestamp 1751266522
transform -1 0 3668 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_146
timestamp 1751266522
transform -1 0 3700 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_373
timestamp 1751266522
transform -1 0 3732 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_374
timestamp 1751266522
transform -1 0 3764 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_464
timestamp 1751266522
transform 1 0 3764 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_14
timestamp 1751266522
transform -1 0 3828 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_372
timestamp 1751266522
transform -1 0 3860 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_66
timestamp 1751266522
transform -1 0 3900 0 -1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_447
timestamp 1751266522
transform -1 0 3932 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_448
timestamp 1751266522
transform 1 0 3932 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_7_0
timestamp 1751266522
transform -1 0 3972 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_7_1
timestamp 1751266522
transform -1 0 3980 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_147
timestamp 1751266522
transform -1 0 4012 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_454
timestamp 1751266522
transform 1 0 4012 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1751266522
transform -1 0 4076 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_64
timestamp 1751266522
transform -1 0 4116 0 -1 305
box -2 -3 42 103
use DFFSR  DFFSR_180
timestamp 1751266522
transform 1 0 4116 0 -1 305
box -2 -3 178 103
use CLKBUF1  CLKBUF1_1
timestamp 1751266522
transform 1 0 4292 0 -1 305
box -2 -3 74 103
use FILL  FILL_3_1
timestamp 1751266522
transform -1 0 4372 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1751266522
transform -1 0 4380 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_3
timestamp 1751266522
transform -1 0 4388 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_4
timestamp 1751266522
transform -1 0 4396 0 -1 305
box -2 -3 10 103
use BUFX2  BUFX2_58
timestamp 1751266522
transform -1 0 28 0 1 305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_46
timestamp 1751266522
transform 1 0 28 0 1 305
box -2 -3 74 103
use DFFSR  DFFSR_87
timestamp 1751266522
transform -1 0 276 0 1 305
box -2 -3 178 103
use BUFX4  BUFX4_214
timestamp 1751266522
transform -1 0 308 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1751266522
transform 1 0 308 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1751266522
transform 1 0 316 0 1 305
box -2 -3 10 103
use DFFSR  DFFSR_27
timestamp 1751266522
transform 1 0 324 0 1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_152
timestamp 1751266522
transform -1 0 532 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_33
timestamp 1751266522
transform -1 0 556 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_156
timestamp 1751266522
transform -1 0 588 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1751266522
transform 1 0 588 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_34
timestamp 1751266522
transform 1 0 620 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_211
timestamp 1751266522
transform 1 0 644 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_102
timestamp 1751266522
transform 1 0 676 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_22
timestamp 1751266522
transform -1 0 884 0 1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_6
timestamp 1751266522
transform 1 0 884 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1751266522
transform 1 0 916 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1751266522
transform 1 0 924 0 1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_5
timestamp 1751266522
transform 1 0 932 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_5
timestamp 1751266522
transform 1 0 964 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1751266522
transform 1 0 996 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_94
timestamp 1751266522
transform 1 0 1020 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1751266522
transform 1 0 1052 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1751266522
transform -1 0 1116 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1751266522
transform 1 0 1116 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_93
timestamp 1751266522
transform 1 0 1148 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1751266522
transform 1 0 1180 0 1 305
box -2 -3 34 103
use INVX1  INVX1_12
timestamp 1751266522
transform -1 0 1228 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_23
timestamp 1751266522
transform 1 0 1228 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_14
timestamp 1751266522
transform 1 0 1260 0 1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_78
timestamp 1751266522
transform -1 0 1332 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1751266522
transform 1 0 1332 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_67
timestamp 1751266522
transform 1 0 1356 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_29
timestamp 1751266522
transform -1 0 1436 0 1 305
box -2 -3 50 103
use FILL  FILL_3_2_0
timestamp 1751266522
transform 1 0 1436 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1751266522
transform 1 0 1444 0 1 305
box -2 -3 10 103
use AOI22X1  AOI22X1_16
timestamp 1751266522
transform 1 0 1452 0 1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_79
timestamp 1751266522
transform -1 0 1524 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1751266522
transform 1 0 1524 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_161
timestamp 1751266522
transform -1 0 1588 0 1 305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_6
timestamp 1751266522
transform 1 0 1588 0 1 305
box -2 -3 74 103
use DFFSR  DFFSR_137
timestamp 1751266522
transform -1 0 1836 0 1 305
box -2 -3 178 103
use AOI22X1  AOI22X1_15
timestamp 1751266522
transform -1 0 1876 0 1 305
box -2 -3 42 103
use CLKBUF1  CLKBUF1_15
timestamp 1751266522
transform -1 0 1948 0 1 305
box -2 -3 74 103
use FILL  FILL_3_3_0
timestamp 1751266522
transform -1 0 1956 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1751266522
transform -1 0 1964 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_234
timestamp 1751266522
transform -1 0 1988 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_626
timestamp 1751266522
transform -1 0 2020 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_178
timestamp 1751266522
transform -1 0 2196 0 1 305
box -2 -3 178 103
use AND2X2  AND2X2_24
timestamp 1751266522
transform 1 0 2196 0 1 305
box -2 -3 34 103
use INVX1  INVX1_114
timestamp 1751266522
transform 1 0 2228 0 1 305
box -2 -3 18 103
use OAI22X1  OAI22X1_110
timestamp 1751266522
transform 1 0 2244 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_538
timestamp 1751266522
transform -1 0 2316 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_537
timestamp 1751266522
transform -1 0 2348 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_536
timestamp 1751266522
transform -1 0 2380 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_176
timestamp 1751266522
transform -1 0 2412 0 1 305
box -2 -3 34 103
use AND2X2  AND2X2_20
timestamp 1751266522
transform -1 0 2444 0 1 305
box -2 -3 34 103
use FILL  FILL_3_4_0
timestamp 1751266522
transform 1 0 2444 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1751266522
transform 1 0 2452 0 1 305
box -2 -3 10 103
use OAI22X1  OAI22X1_102
timestamp 1751266522
transform 1 0 2460 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_509
timestamp 1751266522
transform -1 0 2532 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_508
timestamp 1751266522
transform -1 0 2564 0 1 305
box -2 -3 34 103
use INVX2  INVX2_110
timestamp 1751266522
transform 1 0 2564 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_214
timestamp 1751266522
transform -1 0 2604 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_164
timestamp 1751266522
transform -1 0 2636 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_507
timestamp 1751266522
transform -1 0 2668 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_172
timestamp 1751266522
transform -1 0 2700 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_527
timestamp 1751266522
transform -1 0 2732 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_257
timestamp 1751266522
transform 1 0 2732 0 1 305
box -2 -3 26 103
use DFFSR  DFFSR_151
timestamp 1751266522
transform -1 0 2932 0 1 305
box -2 -3 178 103
use INVX1  INVX1_98
timestamp 1751266522
transform -1 0 2948 0 1 305
box -2 -3 18 103
use FILL  FILL_3_5_0
timestamp 1751266522
transform 1 0 2948 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1751266522
transform 1 0 2956 0 1 305
box -2 -3 10 103
use INVX2  INVX2_111
timestamp 1751266522
transform 1 0 2964 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_439
timestamp 1751266522
transform -1 0 3012 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_62
timestamp 1751266522
transform 1 0 3012 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_440
timestamp 1751266522
transform 1 0 3052 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_243
timestamp 1751266522
transform -1 0 3260 0 1 305
box -2 -3 178 103
use INVX2  INVX2_105
timestamp 1751266522
transform 1 0 3260 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_411
timestamp 1751266522
transform -1 0 3308 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_412
timestamp 1751266522
transform 1 0 3308 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_61
timestamp 1751266522
transform 1 0 3340 0 1 305
box -2 -3 42 103
use BUFX4  BUFX4_12
timestamp 1751266522
transform 1 0 3380 0 1 305
box -2 -3 34 103
use FILL  FILL_3_6_0
timestamp 1751266522
transform -1 0 3420 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1751266522
transform -1 0 3428 0 1 305
box -2 -3 10 103
use DFFSR  DFFSR_226
timestamp 1751266522
transform -1 0 3604 0 1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_506
timestamp 1751266522
transform 1 0 3604 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_266
timestamp 1751266522
transform -1 0 3668 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_172
timestamp 1751266522
transform -1 0 3692 0 1 305
box -2 -3 26 103
use INVX1  INVX1_137
timestamp 1751266522
transform -1 0 3708 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_102
timestamp 1751266522
transform 1 0 3708 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_103
timestamp 1751266522
transform 1 0 3740 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_143
timestamp 1751266522
transform 1 0 3772 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_145
timestamp 1751266522
transform -1 0 3836 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_446
timestamp 1751266522
transform -1 0 3868 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_462
timestamp 1751266522
transform -1 0 3900 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_69
timestamp 1751266522
transform -1 0 3940 0 1 305
box -2 -3 42 103
use AOI22X1  AOI22X1_63
timestamp 1751266522
transform -1 0 3980 0 1 305
box -2 -3 42 103
use FILL  FILL_3_7_0
timestamp 1751266522
transform -1 0 3988 0 1 305
box -2 -3 10 103
use FILL  FILL_3_7_1
timestamp 1751266522
transform -1 0 3996 0 1 305
box -2 -3 10 103
use DFFSR  DFFSR_200
timestamp 1751266522
transform -1 0 4172 0 1 305
box -2 -3 178 103
use NAND3X1  NAND3X1_132
timestamp 1751266522
transform 1 0 4172 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_128
timestamp 1751266522
transform 1 0 4204 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_240
timestamp 1751266522
transform 1 0 4236 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_117
timestamp 1751266522
transform 1 0 4268 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_242
timestamp 1751266522
transform 1 0 4300 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_224
timestamp 1751266522
transform 1 0 4332 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1751266522
transform 1 0 4364 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1751266522
transform 1 0 4372 0 1 305
box -2 -3 10 103
use FILL  FILL_4_3
timestamp 1751266522
transform 1 0 4380 0 1 305
box -2 -3 10 103
use FILL  FILL_4_4
timestamp 1751266522
transform 1 0 4388 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_67
timestamp 1751266522
transform -1 0 28 0 -1 505
box -2 -3 26 103
use DFFSR  DFFSR_96
timestamp 1751266522
transform -1 0 204 0 -1 505
box -2 -3 178 103
use DFFSR  DFFSR_31
timestamp 1751266522
transform 1 0 204 0 -1 505
box -2 -3 178 103
use FILL  FILL_4_0_0
timestamp 1751266522
transform -1 0 388 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1751266522
transform -1 0 396 0 -1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_14
timestamp 1751266522
transform -1 0 468 0 -1 505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_36
timestamp 1751266522
transform 1 0 468 0 -1 505
box -2 -3 74 103
use BUFX2  BUFX2_44
timestamp 1751266522
transform 1 0 540 0 -1 505
box -2 -3 26 103
use DFFSR  DFFSR_20
timestamp 1751266522
transform -1 0 740 0 -1 505
box -2 -3 178 103
use BUFX4  BUFX4_104
timestamp 1751266522
transform 1 0 740 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_95
timestamp 1751266522
transform -1 0 948 0 -1 505
box -2 -3 178 103
use FILL  FILL_4_1_0
timestamp 1751266522
transform -1 0 956 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1751266522
transform -1 0 964 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_3
timestamp 1751266522
transform -1 0 980 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_14
timestamp 1751266522
transform 1 0 980 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1751266522
transform 1 0 1012 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1751266522
transform -1 0 1060 0 -1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_86
timestamp 1751266522
transform -1 0 1092 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_30
timestamp 1751266522
transform 1 0 1092 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_13
timestamp 1751266522
transform 1 0 1132 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1751266522
transform 1 0 1164 0 -1 505
box -2 -3 26 103
use DFFSR  DFFSR_86
timestamp 1751266522
transform 1 0 1188 0 -1 505
box -2 -3 178 103
use BUFX4  BUFX4_116
timestamp 1751266522
transform -1 0 1396 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_604
timestamp 1751266522
transform 1 0 1396 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1751266522
transform 1 0 1428 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1751266522
transform 1 0 1436 0 -1 505
box -2 -3 10 103
use AOI22X1  AOI22X1_29
timestamp 1751266522
transform 1 0 1444 0 -1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_132
timestamp 1751266522
transform 1 0 1484 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_128
timestamp 1751266522
transform -1 0 1532 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_326
timestamp 1751266522
transform 1 0 1532 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_130
timestamp 1751266522
transform 1 0 1564 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_96
timestamp 1751266522
transform -1 0 1612 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_98
timestamp 1751266522
transform -1 0 1636 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_61
timestamp 1751266522
transform 1 0 1636 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_285
timestamp 1751266522
transform -1 0 1684 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_295
timestamp 1751266522
transform 1 0 1684 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_607
timestamp 1751266522
transform -1 0 1748 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_105
timestamp 1751266522
transform 1 0 1748 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_608
timestamp 1751266522
transform 1 0 1764 0 -1 505
box -2 -3 34 103
use AND2X2  AND2X2_22
timestamp 1751266522
transform -1 0 1828 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_605
timestamp 1751266522
transform 1 0 1828 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_226
timestamp 1751266522
transform -1 0 1884 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_3_0
timestamp 1751266522
transform -1 0 1892 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1751266522
transform -1 0 1900 0 -1 505
box -2 -3 10 103
use DFFSR  DFFSR_120
timestamp 1751266522
transform -1 0 2076 0 -1 505
box -2 -3 178 103
use INVX2  INVX2_104
timestamp 1751266522
transform 1 0 2076 0 -1 505
box -2 -3 18 103
use INVX2  INVX2_75
timestamp 1751266522
transform 1 0 2092 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_653
timestamp 1751266522
transform -1 0 2140 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_149
timestamp 1751266522
transform 1 0 2140 0 -1 505
box -2 -3 26 103
use DFFSR  DFFSR_136
timestamp 1751266522
transform -1 0 2340 0 -1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_611
timestamp 1751266522
transform -1 0 2372 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_612
timestamp 1751266522
transform 1 0 2372 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1751266522
transform 1 0 2404 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_4_0
timestamp 1751266522
transform 1 0 2436 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1751266522
transform 1 0 2444 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_16
timestamp 1751266522
transform 1 0 2452 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_689
timestamp 1751266522
transform 1 0 2484 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_74
timestamp 1751266522
transform 1 0 2516 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_217
timestamp 1751266522
transform 1 0 2532 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_258
timestamp 1751266522
transform -1 0 2596 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_171
timestamp 1751266522
transform -1 0 2772 0 -1 505
box -2 -3 178 103
use AOI22X1  AOI22X1_87
timestamp 1751266522
transform 1 0 2772 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_688
timestamp 1751266522
transform 1 0 2812 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_231
timestamp 1751266522
transform -1 0 3020 0 -1 505
box -2 -3 178 103
use FILL  FILL_4_5_0
timestamp 1751266522
transform -1 0 3028 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1751266522
transform -1 0 3036 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_371
timestamp 1751266522
transform -1 0 3068 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_670
timestamp 1751266522
transform -1 0 3100 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_208
timestamp 1751266522
transform -1 0 3132 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_101
timestamp 1751266522
transform 1 0 3132 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_46
timestamp 1751266522
transform 1 0 3164 0 -1 505
box -2 -3 42 103
use BUFX4  BUFX4_157
timestamp 1751266522
transform -1 0 3236 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_438
timestamp 1751266522
transform 1 0 3236 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1751266522
transform -1 0 3300 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_103
timestamp 1751266522
transform -1 0 3316 0 -1 505
box -2 -3 18 103
use DFFSR  DFFSR_242
timestamp 1751266522
transform -1 0 3492 0 -1 505
box -2 -3 178 103
use FILL  FILL_4_6_0
timestamp 1751266522
transform 1 0 3492 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1751266522
transform 1 0 3500 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_81
timestamp 1751266522
transform 1 0 3508 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_36
timestamp 1751266522
transform -1 0 3580 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_370
timestamp 1751266522
transform 1 0 3580 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_100
timestamp 1751266522
transform -1 0 3644 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_381
timestamp 1751266522
transform 1 0 3644 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_380
timestamp 1751266522
transform -1 0 3708 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_121
timestamp 1751266522
transform 1 0 3708 0 -1 505
box -2 -3 18 103
use BUFX4  BUFX4_144
timestamp 1751266522
transform 1 0 3724 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_158
timestamp 1751266522
transform -1 0 3788 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_410
timestamp 1751266522
transform 1 0 3788 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_136
timestamp 1751266522
transform 1 0 3820 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_149
timestamp 1751266522
transform 1 0 3852 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_504
timestamp 1751266522
transform 1 0 3884 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_163
timestamp 1751266522
transform -1 0 3948 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_199
timestamp 1751266522
transform 1 0 3948 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_7_0
timestamp 1751266522
transform -1 0 3988 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_7_1
timestamp 1751266522
transform -1 0 3996 0 -1 505
box -2 -3 10 103
use INVX2  INVX2_138
timestamp 1751266522
transform -1 0 4012 0 -1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_198
timestamp 1751266522
transform 1 0 4012 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_200
timestamp 1751266522
transform -1 0 4076 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_201
timestamp 1751266522
transform 1 0 4076 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_202
timestamp 1751266522
transform -1 0 4140 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_203
timestamp 1751266522
transform -1 0 4172 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1751266522
transform 1 0 4172 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_239
timestamp 1751266522
transform 1 0 4204 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_241
timestamp 1751266522
transform -1 0 4268 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1751266522
transform 1 0 4268 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_244
timestamp 1751266522
transform 1 0 4300 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_243
timestamp 1751266522
transform 1 0 4332 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_221
timestamp 1751266522
transform 1 0 4364 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_17
timestamp 1751266522
transform 1 0 4 0 1 505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_27
timestamp 1751266522
transform 1 0 76 0 1 505
box -2 -3 74 103
use BUFX4  BUFX4_28
timestamp 1751266522
transform 1 0 148 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_213
timestamp 1751266522
transform 1 0 180 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_12
timestamp 1751266522
transform 1 0 212 0 1 505
box -2 -3 178 103
use FILL  FILL_5_0_0
timestamp 1751266522
transform -1 0 396 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1751266522
transform -1 0 404 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_137
timestamp 1751266522
transform -1 0 436 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1751266522
transform 1 0 436 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_42
timestamp 1751266522
transform 1 0 468 0 1 505
box -2 -3 74 103
use BUFX4  BUFX4_195
timestamp 1751266522
transform 1 0 540 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1751266522
transform 1 0 572 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_32
timestamp 1751266522
transform -1 0 780 0 1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_16
timestamp 1751266522
transform 1 0 780 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1751266522
transform -1 0 836 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_98
timestamp 1751266522
transform 1 0 836 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_197
timestamp 1751266522
transform 1 0 868 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1751266522
transform 1 0 900 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1751266522
transform 1 0 908 0 1 505
box -2 -3 10 103
use DFFSR  DFFSR_118
timestamp 1751266522
transform 1 0 916 0 1 505
box -2 -3 178 103
use NAND2X1  NAND2X1_65
timestamp 1751266522
transform -1 0 1116 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_69
timestamp 1751266522
transform -1 0 1148 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_138
timestamp 1751266522
transform 1 0 1148 0 1 505
box -2 -3 178 103
use MUX2X1  MUX2X1_17
timestamp 1751266522
transform 1 0 1324 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_657
timestamp 1751266522
transform 1 0 1372 0 1 505
box -2 -3 34 103
use FILL  FILL_5_2_0
timestamp 1751266522
transform 1 0 1404 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1751266522
transform 1 0 1412 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_603
timestamp 1751266522
transform 1 0 1420 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_134
timestamp 1751266522
transform -1 0 1476 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_324
timestamp 1751266522
transform 1 0 1476 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_329
timestamp 1751266522
transform 1 0 1508 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_131
timestamp 1751266522
transform -1 0 1564 0 1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_76
timestamp 1751266522
transform 1 0 1564 0 1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_283
timestamp 1751266522
transform 1 0 1604 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_327
timestamp 1751266522
transform 1 0 1636 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_294
timestamp 1751266522
transform 1 0 1668 0 1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_64
timestamp 1751266522
transform 1 0 1700 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_106
timestamp 1751266522
transform -1 0 1764 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_104
timestamp 1751266522
transform -1 0 1788 0 1 505
box -2 -3 26 103
use INVX1  INVX1_144
timestamp 1751266522
transform 1 0 1788 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_136
timestamp 1751266522
transform -1 0 1828 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_164
timestamp 1751266522
transform 1 0 1828 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_213
timestamp 1751266522
transform -1 0 1876 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_120
timestamp 1751266522
transform -1 0 1900 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_30
timestamp 1751266522
transform -1 0 1948 0 1 505
box -2 -3 50 103
use FILL  FILL_5_3_0
timestamp 1751266522
transform 1 0 1948 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1751266522
transform 1 0 1956 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_656
timestamp 1751266522
transform 1 0 1964 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_228
timestamp 1751266522
transform -1 0 2020 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_232
timestamp 1751266522
transform 1 0 2020 0 1 505
box -2 -3 26 103
use INVX8  INVX8_24
timestamp 1751266522
transform 1 0 2044 0 1 505
box -2 -3 42 103
use MUX2X1  MUX2X1_42
timestamp 1751266522
transform -1 0 2132 0 1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_241
timestamp 1751266522
transform 1 0 2132 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_625
timestamp 1751266522
transform 1 0 2156 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_225
timestamp 1751266522
transform 1 0 2188 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_618
timestamp 1751266522
transform 1 0 2212 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_652
timestamp 1751266522
transform 1 0 2244 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_241
timestamp 1751266522
transform -1 0 2300 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_239
timestamp 1751266522
transform 1 0 2300 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_223
timestamp 1751266522
transform -1 0 2348 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_23
timestamp 1751266522
transform 1 0 2348 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_610
timestamp 1751266522
transform 1 0 2380 0 1 505
box -2 -3 34 103
use FILL  FILL_5_4_0
timestamp 1751266522
transform -1 0 2420 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1751266522
transform -1 0 2428 0 1 505
box -2 -3 10 103
use DFFSR  DFFSR_150
timestamp 1751266522
transform -1 0 2604 0 1 505
box -2 -3 178 103
use NAND2X1  NAND2X1_215
timestamp 1751266522
transform -1 0 2628 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_252
timestamp 1751266522
transform 1 0 2628 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_17
timestamp 1751266522
transform -1 0 2684 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_240
timestamp 1751266522
transform 1 0 2684 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_213
timestamp 1751266522
transform -1 0 2732 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_260
timestamp 1751266522
transform 1 0 2732 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_18
timestamp 1751266522
transform -1 0 2796 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_251
timestamp 1751266522
transform 1 0 2796 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_216
timestamp 1751266522
transform 1 0 2820 0 1 505
box -2 -3 34 103
use INVX2  INVX2_60
timestamp 1751266522
transform 1 0 2852 0 1 505
box -2 -3 18 103
use FILL  FILL_5_5_0
timestamp 1751266522
transform -1 0 2876 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1751266522
transform -1 0 2884 0 1 505
box -2 -3 10 103
use DFFSR  DFFSR_235
timestamp 1751266522
transform -1 0 3060 0 1 505
box -2 -3 178 103
use INVX2  INVX2_73
timestamp 1751266522
transform 1 0 3060 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_83
timestamp 1751266522
transform 1 0 3076 0 1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_669
timestamp 1751266522
transform 1 0 3116 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_207
timestamp 1751266522
transform -1 0 3180 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_677
timestamp 1751266522
transform 1 0 3180 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_212
timestamp 1751266522
transform 1 0 3212 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_143
timestamp 1751266522
transform 1 0 3244 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_251
timestamp 1751266522
transform -1 0 3308 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_207
timestamp 1751266522
transform 1 0 3308 0 1 505
box -2 -3 26 103
use DFFSR  DFFSR_184
timestamp 1751266522
transform -1 0 3508 0 1 505
box -2 -3 178 103
use FILL  FILL_5_6_0
timestamp 1751266522
transform 1 0 3508 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1751266522
transform 1 0 3516 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_350
timestamp 1751266522
transform 1 0 3524 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_80
timestamp 1751266522
transform -1 0 3588 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_166
timestamp 1751266522
transform -1 0 3612 0 1 505
box -2 -3 26 103
use INVX8  INVX8_17
timestamp 1751266522
transform -1 0 3652 0 1 505
box -2 -3 42 103
use BUFX4  BUFX4_255
timestamp 1751266522
transform 1 0 3652 0 1 505
box -2 -3 34 103
use INVX8  INVX8_14
timestamp 1751266522
transform 1 0 3684 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_171
timestamp 1751266522
transform -1 0 3748 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_254
timestamp 1751266522
transform 1 0 3748 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1751266522
transform -1 0 3804 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_205
timestamp 1751266522
transform -1 0 3828 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_206
timestamp 1751266522
transform -1 0 3852 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_208
timestamp 1751266522
transform 1 0 3852 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_211
timestamp 1751266522
transform 1 0 3876 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_146
timestamp 1751266522
transform 1 0 3900 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_93
timestamp 1751266522
transform 1 0 3932 0 1 505
box -2 -3 34 103
use FILL  FILL_5_7_0
timestamp 1751266522
transform 1 0 3964 0 1 505
box -2 -3 10 103
use FILL  FILL_5_7_1
timestamp 1751266522
transform 1 0 3972 0 1 505
box -2 -3 10 103
use NAND3X1  NAND3X1_162
timestamp 1751266522
transform 1 0 3980 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_92
timestamp 1751266522
transform 1 0 4012 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_161
timestamp 1751266522
transform 1 0 4044 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_118
timestamp 1751266522
transform 1 0 4076 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_177
timestamp 1751266522
transform 1 0 4108 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_131
timestamp 1751266522
transform 1 0 4140 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_133
timestamp 1751266522
transform 1 0 4172 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_129
timestamp 1751266522
transform 1 0 4204 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_119
timestamp 1751266522
transform -1 0 4268 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_114
timestamp 1751266522
transform 1 0 4268 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_225
timestamp 1751266522
transform 1 0 4300 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_226
timestamp 1751266522
transform 1 0 4332 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_223
timestamp 1751266522
transform 1 0 4364 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_38
timestamp 1751266522
transform -1 0 28 0 -1 705
box -2 -3 26 103
use DFFSR  DFFSR_67
timestamp 1751266522
transform -1 0 204 0 -1 705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_38
timestamp 1751266522
transform -1 0 276 0 -1 705
box -2 -3 74 103
use DFFSR  DFFSR_89
timestamp 1751266522
transform -1 0 452 0 -1 705
box -2 -3 178 103
use FILL  FILL_6_0_0
timestamp 1751266522
transform -1 0 460 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1751266522
transform -1 0 468 0 -1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_62
timestamp 1751266522
transform -1 0 540 0 -1 705
box -2 -3 74 103
use DFFSR  DFFSR_73
timestamp 1751266522
transform -1 0 716 0 -1 705
box -2 -3 178 103
use BUFX4  BUFX4_111
timestamp 1751266522
transform 1 0 716 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_109
timestamp 1751266522
transform 1 0 748 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1751266522
transform 1 0 780 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_15
timestamp 1751266522
transform 1 0 796 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1751266522
transform 1 0 828 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_95
timestamp 1751266522
transform 1 0 860 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1751266522
transform 1 0 892 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1751266522
transform 1 0 900 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_105
timestamp 1751266522
transform 1 0 908 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_113
timestamp 1751266522
transform 1 0 940 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_32
timestamp 1751266522
transform 1 0 972 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_87
timestamp 1751266522
transform -1 0 1044 0 -1 705
box -2 -3 34 103
use DFFSR  DFFSR_146
timestamp 1751266522
transform 1 0 1044 0 -1 705
box -2 -3 178 103
use AOI22X1  AOI22X1_8
timestamp 1751266522
transform 1 0 1220 0 -1 705
box -2 -3 42 103
use AOI22X1  AOI22X1_12
timestamp 1751266522
transform 1 0 1260 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_77
timestamp 1751266522
transform -1 0 1332 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1751266522
transform -1 0 1356 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_583
timestamp 1751266522
transform 1 0 1356 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_41
timestamp 1751266522
transform -1 0 1436 0 -1 705
box -2 -3 50 103
use FILL  FILL_6_2_0
timestamp 1751266522
transform 1 0 1436 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1751266522
transform 1 0 1444 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_582
timestamp 1751266522
transform 1 0 1452 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_303
timestamp 1751266522
transform 1 0 1484 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_75
timestamp 1751266522
transform -1 0 1556 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_129
timestamp 1751266522
transform 1 0 1556 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_175
timestamp 1751266522
transform -1 0 1612 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_59
timestamp 1751266522
transform -1 0 1652 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_95
timestamp 1751266522
transform 1 0 1652 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_60
timestamp 1751266522
transform -1 0 1716 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_284
timestamp 1751266522
transform 1 0 1716 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_97
timestamp 1751266522
transform -1 0 1772 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_105
timestamp 1751266522
transform 1 0 1772 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_35
timestamp 1751266522
transform -1 0 1828 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_18
timestamp 1751266522
transform -1 0 1876 0 -1 705
box -2 -3 50 103
use BUFX4  BUFX4_176
timestamp 1751266522
transform -1 0 1908 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_110
timestamp 1751266522
transform 1 0 1908 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_3_0
timestamp 1751266522
transform 1 0 1924 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1751266522
transform 1 0 1932 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_277
timestamp 1751266522
transform 1 0 1940 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_115
timestamp 1751266522
transform 1 0 1972 0 -1 705
box -2 -3 18 103
use DFFSR  DFFSR_169
timestamp 1751266522
transform -1 0 2164 0 -1 705
box -2 -3 178 103
use NOR2X1  NOR2X1_185
timestamp 1751266522
transform -1 0 2188 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_109
timestamp 1751266522
transform 1 0 2188 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_532
timestamp 1751266522
transform -1 0 2260 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_531
timestamp 1751266522
transform -1 0 2292 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_173
timestamp 1751266522
transform -1 0 2324 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_530
timestamp 1751266522
transform 1 0 2324 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_253
timestamp 1751266522
transform 1 0 2356 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_4_0
timestamp 1751266522
transform -1 0 2388 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1751266522
transform -1 0 2396 0 -1 705
box -2 -3 10 103
use DFFSR  DFFSR_148
timestamp 1751266522
transform -1 0 2572 0 -1 705
box -2 -3 178 103
use INVX2  INVX2_125
timestamp 1751266522
transform 1 0 2572 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_223
timestamp 1751266522
transform -1 0 2612 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_188
timestamp 1751266522
transform -1 0 2636 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_196
timestamp 1751266522
transform -1 0 2660 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_698
timestamp 1751266522
transform 1 0 2660 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_651
timestamp 1751266522
transform -1 0 2724 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_80
timestamp 1751266522
transform 1 0 2724 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_222
timestamp 1751266522
transform 1 0 2764 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_574
timestamp 1751266522
transform 1 0 2788 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_199
timestamp 1751266522
transform 1 0 2820 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_198
timestamp 1751266522
transform 1 0 2852 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_159
timestamp 1751266522
transform -1 0 2916 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_126
timestamp 1751266522
transform 1 0 2916 0 -1 705
box -2 -3 18 103
use OAI22X1  OAI22X1_100
timestamp 1751266522
transform 1 0 2932 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_5_0
timestamp 1751266522
transform -1 0 2980 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1751266522
transform -1 0 2988 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_365
timestamp 1751266522
transform -1 0 3020 0 -1 705
box -2 -3 34 103
use DFFSR  DFFSR_182
timestamp 1751266522
transform -1 0 3196 0 -1 705
box -2 -3 178 103
use AOI21X1  AOI21X1_95
timestamp 1751266522
transform -1 0 3228 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_200
timestamp 1751266522
transform -1 0 3252 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_203
timestamp 1751266522
transform -1 0 3276 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_13
timestamp 1751266522
transform -1 0 3308 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_11
timestamp 1751266522
transform -1 0 3340 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1751266522
transform 1 0 3340 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_187
timestamp 1751266522
transform 1 0 3364 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_493
timestamp 1751266522
transform -1 0 3420 0 -1 705
box -2 -3 34 103
use INVX8  INVX8_16
timestamp 1751266522
transform 1 0 3420 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_6_0
timestamp 1751266522
transform 1 0 3460 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1751266522
transform 1 0 3468 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_248
timestamp 1751266522
transform 1 0 3476 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_494
timestamp 1751266522
transform 1 0 3508 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_68
timestamp 1751266522
transform 1 0 3540 0 -1 705
box -2 -3 42 103
use BUFX4  BUFX4_262
timestamp 1751266522
transform -1 0 3612 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_168
timestamp 1751266522
transform -1 0 3636 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_146
timestamp 1751266522
transform -1 0 3652 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_445
timestamp 1751266522
transform -1 0 3684 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_12
timestamp 1751266522
transform 1 0 3684 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1751266522
transform 1 0 3716 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_461
timestamp 1751266522
transform 1 0 3748 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_145
timestamp 1751266522
transform 1 0 3780 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_492
timestamp 1751266522
transform 1 0 3796 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_210
timestamp 1751266522
transform -1 0 3852 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_159
timestamp 1751266522
transform -1 0 3884 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_148
timestamp 1751266522
transform 1 0 3884 0 -1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_207
timestamp 1751266522
transform 1 0 3900 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_174
timestamp 1751266522
transform 1 0 3932 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_7_0
timestamp 1751266522
transform -1 0 3972 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_7_1
timestamp 1751266522
transform -1 0 3980 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_94
timestamp 1751266522
transform -1 0 4012 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_173
timestamp 1751266522
transform 1 0 4012 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_175
timestamp 1751266522
transform -1 0 4076 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_176
timestamp 1751266522
transform 1 0 4076 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_178
timestamp 1751266522
transform -1 0 4140 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1751266522
transform 1 0 4140 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1751266522
transform -1 0 4204 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_130
timestamp 1751266522
transform 1 0 4204 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1751266522
transform -1 0 4268 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_116
timestamp 1751266522
transform 1 0 4268 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_115
timestamp 1751266522
transform 1 0 4300 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_51
timestamp 1751266522
transform 1 0 4332 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1751266522
transform 1 0 4364 0 -1 705
box -2 -3 34 103
use BUFX2  BUFX2_27
timestamp 1751266522
transform -1 0 28 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_55
timestamp 1751266522
transform -1 0 52 0 1 705
box -2 -3 26 103
use DFFSR  DFFSR_84
timestamp 1751266522
transform -1 0 228 0 1 705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_59
timestamp 1751266522
transform 1 0 228 0 1 705
box -2 -3 74 103
use OAI21X1  OAI21X1_150
timestamp 1751266522
transform 1 0 300 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_4
timestamp 1751266522
transform 1 0 332 0 1 705
box -2 -3 74 103
use FILL  FILL_7_0_0
timestamp 1751266522
transform -1 0 412 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1751266522
transform -1 0 420 0 1 705
box -2 -3 10 103
use DFFSR  DFFSR_30
timestamp 1751266522
transform -1 0 596 0 1 705
box -2 -3 178 103
use BUFX4  BUFX4_106
timestamp 1751266522
transform 1 0 596 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_1
timestamp 1751266522
transform -1 0 660 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1751266522
transform 1 0 660 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_12
timestamp 1751266522
transform -1 0 724 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1751266522
transform -1 0 756 0 1 705
box -2 -3 34 103
use INVX1  INVX1_6
timestamp 1751266522
transform -1 0 772 0 1 705
box -2 -3 18 103
use DFFSR  DFFSR_142
timestamp 1751266522
transform 1 0 772 0 1 705
box -2 -3 178 103
use FILL  FILL_7_1_0
timestamp 1751266522
transform 1 0 948 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1751266522
transform 1 0 956 0 1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_35
timestamp 1751266522
transform 1 0 964 0 1 705
box -2 -3 74 103
use NAND2X1  NAND2X1_37
timestamp 1751266522
transform -1 0 1060 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1751266522
transform -1 0 1092 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_70
timestamp 1751266522
transform -1 0 1124 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_5
timestamp 1751266522
transform -1 0 1156 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1751266522
transform -1 0 1180 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_75
timestamp 1751266522
transform -1 0 1212 0 1 705
box -2 -3 34 103
use DFFSR  DFFSR_147
timestamp 1751266522
transform -1 0 1388 0 1 705
box -2 -3 178 103
use INVX1  INVX1_24
timestamp 1751266522
transform -1 0 1404 0 1 705
box -2 -3 18 103
use INVX1  INVX1_25
timestamp 1751266522
transform -1 0 1420 0 1 705
box -2 -3 18 103
use FILL  FILL_7_2_0
timestamp 1751266522
transform -1 0 1428 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1751266522
transform -1 0 1436 0 1 705
box -2 -3 10 103
use INVX1  INVX1_30
timestamp 1751266522
transform -1 0 1452 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1751266522
transform 1 0 1452 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_331
timestamp 1751266522
transform 1 0 1492 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_262
timestamp 1751266522
transform 1 0 1524 0 1 705
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1751266522
transform -1 0 1572 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_328
timestamp 1751266522
transform 1 0 1572 0 1 705
box -2 -3 34 103
use INVX1  INVX1_108
timestamp 1751266522
transform 1 0 1604 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_11
timestamp 1751266522
transform 1 0 1620 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_286
timestamp 1751266522
transform 1 0 1660 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_272
timestamp 1751266522
transform 1 0 1692 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_336
timestamp 1751266522
transform 1 0 1724 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1751266522
transform -1 0 1788 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_315
timestamp 1751266522
transform -1 0 1820 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_138
timestamp 1751266522
transform -1 0 1844 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_222
timestamp 1751266522
transform -1 0 1868 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_214
timestamp 1751266522
transform 1 0 1868 0 1 705
box -2 -3 26 103
use INVX2  INVX2_98
timestamp 1751266522
transform 1 0 1892 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_221
timestamp 1751266522
transform 1 0 1908 0 1 705
box -2 -3 26 103
use FILL  FILL_7_3_0
timestamp 1751266522
transform -1 0 1940 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1751266522
transform -1 0 1948 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_606
timestamp 1751266522
transform -1 0 1980 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_243
timestamp 1751266522
transform -1 0 2004 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_581
timestamp 1751266522
transform 1 0 2004 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_602
timestamp 1751266522
transform 1 0 2036 0 1 705
box -2 -3 34 103
use DFFSR  DFFSR_199
timestamp 1751266522
transform -1 0 2244 0 1 705
box -2 -3 178 103
use BUFX4  BUFX4_273
timestamp 1751266522
transform 1 0 2244 0 1 705
box -2 -3 34 103
use INVX1  INVX1_118
timestamp 1751266522
transform 1 0 2276 0 1 705
box -2 -3 18 103
use AND2X2  AND2X2_19
timestamp 1751266522
transform 1 0 2292 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_151
timestamp 1751266522
transform -1 0 2356 0 1 705
box -2 -3 34 103
use INVX2  INVX2_149
timestamp 1751266522
transform 1 0 2356 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_81
timestamp 1751266522
transform 1 0 2372 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_579
timestamp 1751266522
transform 1 0 2412 0 1 705
box -2 -3 34 103
use FILL  FILL_7_4_0
timestamp 1751266522
transform 1 0 2444 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1751266522
transform 1 0 2452 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_202
timestamp 1751266522
transform 1 0 2460 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1751266522
transform -1 0 2524 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_200
timestamp 1751266522
transform 1 0 2524 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_204
timestamp 1751266522
transform 1 0 2556 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_221
timestamp 1751266522
transform -1 0 2604 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_197
timestamp 1751266522
transform -1 0 2636 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_572
timestamp 1751266522
transform -1 0 2668 0 1 705
box -2 -3 34 103
use DFFSR  DFFSR_201
timestamp 1751266522
transform -1 0 2844 0 1 705
box -2 -3 178 103
use AOI22X1  AOI22X1_79
timestamp 1751266522
transform -1 0 2884 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_499
timestamp 1751266522
transform -1 0 2916 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_500
timestamp 1751266522
transform 1 0 2916 0 1 705
box -2 -3 34 103
use FILL  FILL_7_5_0
timestamp 1751266522
transform 1 0 2948 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1751266522
transform 1 0 2956 0 1 705
box -2 -3 10 103
use INVX2  INVX2_109
timestamp 1751266522
transform 1 0 2964 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_498
timestamp 1751266522
transform -1 0 3012 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_161
timestamp 1751266522
transform -1 0 3044 0 1 705
box -2 -3 34 103
use DFFSR  DFFSR_216
timestamp 1751266522
transform -1 0 3220 0 1 705
box -2 -3 178 103
use NOR2X1  NOR2X1_183
timestamp 1751266522
transform -1 0 3244 0 1 705
box -2 -3 26 103
use INVX2  INVX2_133
timestamp 1751266522
transform 1 0 3244 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_56
timestamp 1751266522
transform 1 0 3260 0 1 705
box -2 -3 42 103
use INVX2  INVX2_135
timestamp 1751266522
transform 1 0 3300 0 1 705
box -2 -3 18 103
use DFFSR  DFFSR_214
timestamp 1751266522
transform -1 0 3492 0 1 705
box -2 -3 178 103
use FILL  FILL_7_6_0
timestamp 1751266522
transform 1 0 3492 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1751266522
transform 1 0 3500 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_399
timestamp 1751266522
transform 1 0 3508 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_126
timestamp 1751266522
transform -1 0 3572 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1751266522
transform 1 0 3572 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_505
timestamp 1751266522
transform -1 0 3628 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1751266522
transform 1 0 3628 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_54
timestamp 1751266522
transform 1 0 3660 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_148
timestamp 1751266522
transform -1 0 3716 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_409
timestamp 1751266522
transform 1 0 3716 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_155
timestamp 1751266522
transform 1 0 3748 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1751266522
transform 1 0 3780 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_208
timestamp 1751266522
transform 1 0 3804 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_165
timestamp 1751266522
transform 1 0 3836 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_209
timestamp 1751266522
transform -1 0 3900 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_148
timestamp 1751266522
transform 1 0 3900 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_164
timestamp 1751266522
transform 1 0 3932 0 1 705
box -2 -3 34 103
use FILL  FILL_7_7_0
timestamp 1751266522
transform 1 0 3964 0 1 705
box -2 -3 10 103
use FILL  FILL_7_7_1
timestamp 1751266522
transform 1 0 3972 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_144
timestamp 1751266522
transform 1 0 3980 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_205
timestamp 1751266522
transform 1 0 4012 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_163
timestamp 1751266522
transform -1 0 4076 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_73
timestamp 1751266522
transform -1 0 4108 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_218
timestamp 1751266522
transform 1 0 4108 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_56
timestamp 1751266522
transform -1 0 4172 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_134
timestamp 1751266522
transform -1 0 4204 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_219
timestamp 1751266522
transform 1 0 4204 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_71
timestamp 1751266522
transform 1 0 4236 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_61
timestamp 1751266522
transform -1 0 4300 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_215
timestamp 1751266522
transform 1 0 4300 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_141
timestamp 1751266522
transform -1 0 4364 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_140
timestamp 1751266522
transform -1 0 4396 0 1 705
box -2 -3 34 103
use BUFX2  BUFX2_42
timestamp 1751266522
transform -1 0 28 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_5
timestamp 1751266522
transform -1 0 52 0 -1 905
box -2 -3 26 103
use DFFSR  DFFSR_71
timestamp 1751266522
transform -1 0 228 0 -1 905
box -2 -3 178 103
use OAI21X1  OAI21X1_128
timestamp 1751266522
transform 1 0 228 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_32
timestamp 1751266522
transform -1 0 332 0 -1 905
box -2 -3 74 103
use FILL  FILL_8_0_0
timestamp 1751266522
transform -1 0 340 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1751266522
transform -1 0 348 0 -1 905
box -2 -3 10 103
use DFFSR  DFFSR_25
timestamp 1751266522
transform -1 0 524 0 -1 905
box -2 -3 178 103
use BUFX4  BUFX4_120
timestamp 1751266522
transform -1 0 556 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_11
timestamp 1751266522
transform 1 0 556 0 -1 905
box -2 -3 74 103
use BUFX4  BUFX4_112
timestamp 1751266522
transform 1 0 628 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1751266522
transform 1 0 660 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1751266522
transform 1 0 692 0 -1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_3
timestamp 1751266522
transform 1 0 708 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_1
timestamp 1751266522
transform 1 0 740 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_108
timestamp 1751266522
transform 1 0 772 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1751266522
transform 1 0 804 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1751266522
transform 1 0 828 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1751266522
transform 1 0 836 0 -1 905
box -2 -3 10 103
use DFFSR  DFFSR_122
timestamp 1751266522
transform 1 0 844 0 -1 905
box -2 -3 178 103
use NOR2X1  NOR2X1_4
timestamp 1751266522
transform 1 0 1020 0 -1 905
box -2 -3 26 103
use DFFSR  DFFSR_123
timestamp 1751266522
transform -1 0 1220 0 -1 905
box -2 -3 178 103
use NAND2X1  NAND2X1_27
timestamp 1751266522
transform 1 0 1220 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_54
timestamp 1751266522
transform -1 0 1268 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_29
timestamp 1751266522
transform 1 0 1268 0 -1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_13
timestamp 1751266522
transform 1 0 1292 0 -1 905
box -2 -3 42 103
use INVX1  INVX1_31
timestamp 1751266522
transform -1 0 1348 0 -1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_7
timestamp 1751266522
transform 1 0 1348 0 -1 905
box -2 -3 42 103
use BUFX4  BUFX4_222
timestamp 1751266522
transform 1 0 1388 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_2_0
timestamp 1751266522
transform 1 0 1420 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1751266522
transform 1 0 1428 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_113
timestamp 1751266522
transform 1 0 1436 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_112
timestamp 1751266522
transform 1 0 1460 0 -1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_67
timestamp 1751266522
transform -1 0 1524 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_304
timestamp 1751266522
transform -1 0 1556 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_325
timestamp 1751266522
transform -1 0 1588 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_292
timestamp 1751266522
transform 1 0 1588 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1751266522
transform -1 0 1652 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_78
timestamp 1751266522
transform 1 0 1652 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_337
timestamp 1751266522
transform 1 0 1676 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_103
timestamp 1751266522
transform -1 0 1732 0 -1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_63
timestamp 1751266522
transform 1 0 1732 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_293
timestamp 1751266522
transform -1 0 1804 0 -1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_80
timestamp 1751266522
transform 1 0 1804 0 -1 905
box -2 -3 42 103
use BUFX4  BUFX4_221
timestamp 1751266522
transform -1 0 1876 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_3_0
timestamp 1751266522
transform -1 0 1884 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1751266522
transform -1 0 1892 0 -1 905
box -2 -3 10 103
use DFFSR  DFFSR_152
timestamp 1751266522
transform -1 0 2068 0 -1 905
box -2 -3 178 103
use NOR2X1  NOR2X1_237
timestamp 1751266522
transform -1 0 2092 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_230
timestamp 1751266522
transform -1 0 2116 0 -1 905
box -2 -3 26 103
use DFFSR  DFFSR_154
timestamp 1751266522
transform -1 0 2292 0 -1 905
box -2 -3 178 103
use INVX2  INVX2_134
timestamp 1751266522
transform 1 0 2292 0 -1 905
box -2 -3 18 103
use BUFX4  BUFX4_127
timestamp 1751266522
transform 1 0 2308 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_200
timestamp 1751266522
transform -1 0 2364 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_228
timestamp 1751266522
transform 1 0 2364 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_613
timestamp 1751266522
transform -1 0 2420 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_216
timestamp 1751266522
transform 1 0 2420 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_4_0
timestamp 1751266522
transform 1 0 2444 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1751266522
transform 1 0 2452 0 -1 905
box -2 -3 10 103
use AOI22X1  AOI22X1_78
timestamp 1751266522
transform 1 0 2460 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_570
timestamp 1751266522
transform 1 0 2500 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_195
timestamp 1751266522
transform -1 0 2564 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1751266522
transform -1 0 2588 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_196
timestamp 1751266522
transform -1 0 2620 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_571
timestamp 1751266522
transform 1 0 2620 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_218
timestamp 1751266522
transform -1 0 2676 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_203
timestamp 1751266522
transform -1 0 2708 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_256
timestamp 1751266522
transform -1 0 2740 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_252
timestamp 1751266522
transform -1 0 2764 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_65
timestamp 1751266522
transform 1 0 2764 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_580
timestamp 1751266522
transform -1 0 2812 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_99
timestamp 1751266522
transform 1 0 2812 0 -1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_89
timestamp 1751266522
transform -1 0 2868 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_444
timestamp 1751266522
transform -1 0 2900 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_443
timestamp 1751266522
transform -1 0 2932 0 -1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_90
timestamp 1751266522
transform -1 0 2972 0 -1 905
box -2 -3 42 103
use FILL  FILL_8_5_0
timestamp 1751266522
transform -1 0 2980 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1751266522
transform -1 0 2988 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_452
timestamp 1751266522
transform -1 0 3020 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_451
timestamp 1751266522
transform -1 0 3052 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_367
timestamp 1751266522
transform -1 0 3084 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_155
timestamp 1751266522
transform -1 0 3100 0 -1 905
box -2 -3 18 103
use INVX2  INVX2_97
timestamp 1751266522
transform 1 0 3100 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_250
timestamp 1751266522
transform 1 0 3116 0 -1 905
box -2 -3 26 103
use INVX8  INVX8_19
timestamp 1751266522
transform 1 0 3140 0 -1 905
box -2 -3 42 103
use AOI22X1  AOI22X1_43
timestamp 1751266522
transform 1 0 3180 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_533
timestamp 1751266522
transform -1 0 3252 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_400
timestamp 1751266522
transform 1 0 3252 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_127
timestamp 1751266522
transform 1 0 3284 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_404
timestamp 1751266522
transform -1 0 3348 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_364
timestamp 1751266522
transform 1 0 3348 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_94
timestamp 1751266522
transform -1 0 3412 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_131
timestamp 1751266522
transform 1 0 3412 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_58
timestamp 1751266522
transform 1 0 3444 0 -1 905
box -2 -3 42 103
use FILL  FILL_8_6_0
timestamp 1751266522
transform -1 0 3492 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1751266522
transform -1 0 3500 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_408
timestamp 1751266522
transform -1 0 3532 0 -1 905
box -2 -3 34 103
use DFFSR  DFFSR_212
timestamp 1751266522
transform -1 0 3708 0 -1 905
box -2 -3 178 103
use AOI21X1  AOI21X1_135
timestamp 1751266522
transform 1 0 3708 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_403
timestamp 1751266522
transform -1 0 3772 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_60
timestamp 1751266522
transform 1 0 3772 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_407
timestamp 1751266522
transform 1 0 3812 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_134
timestamp 1751266522
transform -1 0 3876 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_203
timestamp 1751266522
transform -1 0 3900 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_209
timestamp 1751266522
transform 1 0 3900 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_147
timestamp 1751266522
transform 1 0 3924 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_166
timestamp 1751266522
transform -1 0 3988 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_7_0
timestamp 1751266522
transform 1 0 3988 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_7_1
timestamp 1751266522
transform 1 0 3996 0 -1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_143
timestamp 1751266522
transform 1 0 4004 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_145
timestamp 1751266522
transform -1 0 4068 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_204
timestamp 1751266522
transform 1 0 4068 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_206
timestamp 1751266522
transform -1 0 4132 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_44
timestamp 1751266522
transform 1 0 4132 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_51
timestamp 1751266522
transform 1 0 4164 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_150
timestamp 1751266522
transform -1 0 4212 0 -1 905
box -2 -3 18 103
use BUFX4  BUFX4_60
timestamp 1751266522
transform -1 0 4244 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_72
timestamp 1751266522
transform -1 0 4276 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_220
timestamp 1751266522
transform -1 0 4308 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_216
timestamp 1751266522
transform 1 0 4308 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_217
timestamp 1751266522
transform -1 0 4372 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1751266522
transform -1 0 4380 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1751266522
transform -1 0 4388 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_3
timestamp 1751266522
transform -1 0 4396 0 -1 905
box -2 -3 10 103
use BUFX2  BUFX2_17
timestamp 1751266522
transform -1 0 28 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_43
timestamp 1751266522
transform -1 0 52 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_72
timestamp 1751266522
transform -1 0 228 0 1 905
box -2 -3 178 103
use OAI21X1  OAI21X1_140
timestamp 1751266522
transform 1 0 228 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_63
timestamp 1751266522
transform -1 0 284 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_15
timestamp 1751266522
transform -1 0 460 0 1 905
box -2 -3 178 103
use FILL  FILL_9_0_0
timestamp 1751266522
transform -1 0 468 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1751266522
transform -1 0 476 0 1 905
box -2 -3 10 103
use DFFSR  DFFSR_92
timestamp 1751266522
transform -1 0 652 0 1 905
box -2 -3 178 103
use INVX2  INVX2_12
timestamp 1751266522
transform 1 0 652 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_54
timestamp 1751266522
transform 1 0 668 0 1 905
box -2 -3 34 103
use DFFSR  DFFSR_3
timestamp 1751266522
transform -1 0 876 0 1 905
box -2 -3 178 103
use BUFX4  BUFX4_110
timestamp 1751266522
transform -1 0 908 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1751266522
transform 1 0 908 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1751266522
transform 1 0 916 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_107
timestamp 1751266522
transform 1 0 924 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1751266522
transform 1 0 956 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_41
timestamp 1751266522
transform -1 0 1004 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_8
timestamp 1751266522
transform 1 0 1004 0 1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_18
timestamp 1751266522
transform 1 0 1028 0 1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_7
timestamp 1751266522
transform 1 0 1068 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_35
timestamp 1751266522
transform -1 0 1148 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_648
timestamp 1751266522
transform 1 0 1148 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1751266522
transform -1 0 1228 0 1 905
box -2 -3 50 103
use BUFX4  BUFX4_124
timestamp 1751266522
transform -1 0 1260 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_702
timestamp 1751266522
transform 1 0 1260 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_596
timestamp 1751266522
transform 1 0 1292 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_685
timestamp 1751266522
transform -1 0 1356 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_45
timestamp 1751266522
transform 1 0 1356 0 1 905
box -2 -3 50 103
use INVX1  INVX1_28
timestamp 1751266522
transform -1 0 1420 0 1 905
box -2 -3 18 103
use FILL  FILL_9_2_0
timestamp 1751266522
transform 1 0 1420 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1751266522
transform 1 0 1428 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_701
timestamp 1751266522
transform 1 0 1436 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_647
timestamp 1751266522
transform 1 0 1468 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_172
timestamp 1751266522
transform -1 0 1532 0 1 905
box -2 -3 34 103
use INVX1  INVX1_26
timestamp 1751266522
transform -1 0 1548 0 1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_1
timestamp 1751266522
transform 1 0 1548 0 1 905
box -2 -3 42 103
use INVX1  INVX1_32
timestamp 1751266522
transform -1 0 1604 0 1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_77
timestamp 1751266522
transform -1 0 1644 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_133
timestamp 1751266522
transform 1 0 1644 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_79
timestamp 1751266522
transform -1 0 1700 0 1 905
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1751266522
transform -1 0 1716 0 1 905
box -2 -3 18 103
use INVX1  INVX1_111
timestamp 1751266522
transform 1 0 1716 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_39
timestamp 1751266522
transform -1 0 1764 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_80
timestamp 1751266522
transform -1 0 1796 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_296
timestamp 1751266522
transform 1 0 1796 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_139
timestamp 1751266522
transform 1 0 1828 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_334
timestamp 1751266522
transform -1 0 1884 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_313
timestamp 1751266522
transform -1 0 1916 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_122
timestamp 1751266522
transform 1 0 1916 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1751266522
transform 1 0 1940 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1751266522
transform 1 0 1948 0 1 905
box -2 -3 10 103
use INVX1  INVX1_123
timestamp 1751266522
transform 1 0 1956 0 1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_44
timestamp 1751266522
transform 1 0 1972 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_36
timestamp 1751266522
transform -1 0 2068 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_48
timestamp 1751266522
transform -1 0 2116 0 1 905
box -2 -3 50 103
use INVX2  INVX2_113
timestamp 1751266522
transform 1 0 2116 0 1 905
box -2 -3 18 103
use INVX2  INVX2_107
timestamp 1751266522
transform 1 0 2132 0 1 905
box -2 -3 18 103
use DFFSR  DFFSR_162
timestamp 1751266522
transform -1 0 2324 0 1 905
box -2 -3 178 103
use AOI22X1  AOI22X1_74
timestamp 1751266522
transform 1 0 2324 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_173
timestamp 1751266522
transform -1 0 2388 0 1 905
box -2 -3 26 103
use INVX1  INVX1_94
timestamp 1751266522
transform 1 0 2388 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_7
timestamp 1751266522
transform -1 0 2436 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1751266522
transform 1 0 2436 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1751266522
transform 1 0 2444 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_547
timestamp 1751266522
transform 1 0 2452 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_182
timestamp 1751266522
transform 1 0 2484 0 1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_76
timestamp 1751266522
transform 1 0 2516 0 1 905
box -2 -3 42 103
use INVX8  INVX8_23
timestamp 1751266522
transform -1 0 2596 0 1 905
box -2 -3 42 103
use INVX2  INVX2_62
timestamp 1751266522
transform 1 0 2596 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_566
timestamp 1751266522
transform 1 0 2612 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_191
timestamp 1751266522
transform -1 0 2676 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_690
timestamp 1751266522
transform 1 0 2676 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_218
timestamp 1751266522
transform -1 0 2740 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_198
timestamp 1751266522
transform 1 0 2740 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_573
timestamp 1751266522
transform 1 0 2764 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1751266522
transform 1 0 2796 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_442
timestamp 1751266522
transform 1 0 2828 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_450
timestamp 1751266522
transform -1 0 2892 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_146
timestamp 1751266522
transform 1 0 2892 0 1 905
box -2 -3 34 103
use FILL  FILL_9_5_0
timestamp 1751266522
transform -1 0 2932 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1751266522
transform -1 0 2940 0 1 905
box -2 -3 10 103
use DFFSR  DFFSR_234
timestamp 1751266522
transform -1 0 3116 0 1 905
box -2 -3 178 103
use OAI21X1  OAI21X1_402
timestamp 1751266522
transform -1 0 3148 0 1 905
box -2 -3 34 103
use INVX2  INVX2_64
timestamp 1751266522
transform 1 0 3148 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_246
timestamp 1751266522
transform -1 0 3188 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_215
timestamp 1751266522
transform -1 0 3364 0 1 905
box -2 -3 178 103
use INVX2  INVX2_124
timestamp 1751266522
transform 1 0 3364 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_162
timestamp 1751266522
transform -1 0 3404 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_129
timestamp 1751266522
transform 1 0 3404 0 1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_57
timestamp 1751266522
transform 1 0 3436 0 1 905
box -2 -3 42 103
use FILL  FILL_9_6_0
timestamp 1751266522
transform -1 0 3484 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1751266522
transform -1 0 3492 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_389
timestamp 1751266522
transform -1 0 3524 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_245
timestamp 1751266522
transform 1 0 3524 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_197
timestamp 1751266522
transform 1 0 3556 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_401
timestamp 1751266522
transform 1 0 3580 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_128
timestamp 1751266522
transform 1 0 3612 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_126
timestamp 1751266522
transform 1 0 3644 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_261
timestamp 1751266522
transform -1 0 3708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_467
timestamp 1751266522
transform 1 0 3708 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_130
timestamp 1751266522
transform -1 0 3772 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1751266522
transform 1 0 3772 0 1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_67
timestamp 1751266522
transform 1 0 3796 0 1 905
box -2 -3 42 103
use CLKBUF1  CLKBUF1_16
timestamp 1751266522
transform -1 0 3908 0 1 905
box -2 -3 74 103
use OAI21X1  OAI21X1_465
timestamp 1751266522
transform 1 0 3908 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_150
timestamp 1751266522
transform -1 0 3972 0 1 905
box -2 -3 34 103
use FILL  FILL_9_7_0
timestamp 1751266522
transform 1 0 3972 0 1 905
box -2 -3 10 103
use FILL  FILL_9_7_1
timestamp 1751266522
transform 1 0 3980 0 1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_96
timestamp 1751266522
transform 1 0 3988 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_101
timestamp 1751266522
transform 1 0 4020 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_103
timestamp 1751266522
transform -1 0 4084 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_149
timestamp 1751266522
transform 1 0 4084 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_246
timestamp 1751266522
transform 1 0 4116 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_206
timestamp 1751266522
transform -1 0 4180 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_249
timestamp 1751266522
transform 1 0 4180 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_248
timestamp 1751266522
transform 1 0 4212 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_182
timestamp 1751266522
transform 1 0 4244 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1751266522
transform 1 0 4276 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_62
timestamp 1751266522
transform 1 0 4308 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1751266522
transform -1 0 4372 0 1 905
box -2 -3 34 103
use FILL  FILL_10_1
timestamp 1751266522
transform 1 0 4372 0 1 905
box -2 -3 10 103
use FILL  FILL_10_2
timestamp 1751266522
transform 1 0 4380 0 1 905
box -2 -3 10 103
use FILL  FILL_10_3
timestamp 1751266522
transform 1 0 4388 0 1 905
box -2 -3 10 103
use BUFX2  BUFX2_12
timestamp 1751266522
transform -1 0 28 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_62
timestamp 1751266522
transform -1 0 52 0 -1 1105
box -2 -3 26 103
use DFFSR  DFFSR_91
timestamp 1751266522
transform -1 0 228 0 -1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_135
timestamp 1751266522
transform 1 0 228 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_10
timestamp 1751266522
transform -1 0 436 0 -1 1105
box -2 -3 178 103
use FILL  FILL_10_0_0
timestamp 1751266522
transform 1 0 436 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1751266522
transform 1 0 444 0 -1 1105
box -2 -3 10 103
use DFFSR  DFFSR_5
timestamp 1751266522
transform 1 0 452 0 -1 1105
box -2 -3 178 103
use INVX2  INVX2_14
timestamp 1751266522
transform 1 0 628 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_58
timestamp 1751266522
transform 1 0 644 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_29
timestamp 1751266522
transform 1 0 676 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1751266522
transform 1 0 708 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_57
timestamp 1751266522
transform 1 0 740 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_140
timestamp 1751266522
transform 1 0 772 0 -1 1105
box -2 -3 178 103
use FILL  FILL_10_1_0
timestamp 1751266522
transform 1 0 948 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1751266522
transform 1 0 956 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_8
timestamp 1751266522
transform 1 0 964 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_15
timestamp 1751266522
transform -1 0 1020 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_22
timestamp 1751266522
transform 1 0 1020 0 -1 1105
box -2 -3 42 103
use NAND3X1  NAND3X1_80
timestamp 1751266522
transform 1 0 1060 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_145
timestamp 1751266522
transform 1 0 1092 0 -1 1105
box -2 -3 178 103
use MUX2X1  MUX2X1_23
timestamp 1751266522
transform 1 0 1268 0 -1 1105
box -2 -3 50 103
use OAI22X1  OAI22X1_19
timestamp 1751266522
transform 1 0 1316 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_157
timestamp 1751266522
transform -1 0 1380 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_37
timestamp 1751266522
transform -1 0 1396 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_36
timestamp 1751266522
transform -1 0 1412 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_2_0
timestamp 1751266522
transform 1 0 1412 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1751266522
transform 1 0 1420 0 -1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_43
timestamp 1751266522
transform 1 0 1428 0 -1 1105
box -2 -3 50 103
use OAI22X1  OAI22X1_78
timestamp 1751266522
transform 1 0 1476 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_135
timestamp 1751266522
transform -1 0 1540 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_662
timestamp 1751266522
transform 1 0 1540 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_661
timestamp 1751266522
transform 1 0 1572 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_144
timestamp 1751266522
transform 1 0 1604 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_333
timestamp 1751266522
transform 1 0 1628 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_330
timestamp 1751266522
transform -1 0 1692 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_259
timestamp 1751266522
transform 1 0 1692 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_224
timestamp 1751266522
transform -1 0 1756 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_137
timestamp 1751266522
transform 1 0 1756 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_79
timestamp 1751266522
transform 1 0 1780 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_338
timestamp 1751266522
transform 1 0 1820 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_121
timestamp 1751266522
transform 1 0 1852 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_71
timestamp 1751266522
transform 1 0 1876 0 -1 1105
box -2 -3 42 103
use FILL  FILL_10_3_0
timestamp 1751266522
transform 1 0 1916 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1751266522
transform 1 0 1924 0 -1 1105
box -2 -3 10 103
use OAI22X1  OAI22X1_72
timestamp 1751266522
transform 1 0 1932 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_123
timestamp 1751266522
transform 1 0 1972 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_317
timestamp 1751266522
transform 1 0 1996 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_99
timestamp 1751266522
transform 1 0 2028 0 -1 1105
box -2 -3 18 103
use BUFX4  BUFX4_179
timestamp 1751266522
transform 1 0 2044 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_229
timestamp 1751266522
transform -1 0 2100 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_615
timestamp 1751266522
transform -1 0 2132 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_138
timestamp 1751266522
transform 1 0 2132 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_204
timestamp 1751266522
transform -1 0 2172 0 -1 1105
box -2 -3 26 103
use DFFSR  DFFSR_135
timestamp 1751266522
transform -1 0 2348 0 -1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_616
timestamp 1751266522
transform 1 0 2348 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_206
timestamp 1751266522
transform 1 0 2380 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_161
timestamp 1751266522
transform -1 0 2428 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_4_0
timestamp 1751266522
transform 1 0 2428 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1751266522
transform 1 0 2436 0 -1 1105
box -2 -3 10 103
use BUFX4  BUFX4_5
timestamp 1751266522
transform 1 0 2444 0 -1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_19
timestamp 1751266522
transform 1 0 2476 0 -1 1105
box -2 -3 74 103
use INVX2  INVX2_77
timestamp 1751266522
transform 1 0 2548 0 -1 1105
box -2 -3 18 103
use BUFX4  BUFX4_259
timestamp 1751266522
transform -1 0 2596 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_257
timestamp 1751266522
transform 1 0 2596 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_88
timestamp 1751266522
transform 1 0 2628 0 -1 1105
box -2 -3 42 103
use DFFSR  DFFSR_155
timestamp 1751266522
transform -1 0 2844 0 -1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_202
timestamp 1751266522
transform 1 0 2844 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_172
timestamp 1751266522
transform -1 0 2892 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_497
timestamp 1751266522
transform -1 0 2924 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_496
timestamp 1751266522
transform -1 0 2956 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_5_0
timestamp 1751266522
transform -1 0 2964 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1751266522
transform -1 0 2972 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_157
timestamp 1751266522
transform -1 0 3004 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_222
timestamp 1751266522
transform -1 0 3180 0 -1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_248
timestamp 1751266522
transform -1 0 3204 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_180
timestamp 1751266522
transform 1 0 3204 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_97
timestamp 1751266522
transform 1 0 3228 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_541
timestamp 1751266522
transform 1 0 3260 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_676
timestamp 1751266522
transform -1 0 3324 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_449
timestamp 1751266522
transform 1 0 3324 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1751266522
transform 1 0 3356 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_147
timestamp 1751266522
transform -1 0 3404 0 -1 1105
box -2 -3 18 103
use BUFX4  BUFX4_53
timestamp 1751266522
transform -1 0 3436 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_457
timestamp 1751266522
transform 1 0 3436 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_6_0
timestamp 1751266522
transform -1 0 3476 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1751266522
transform -1 0 3484 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_390
timestamp 1751266522
transform -1 0 3516 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_148
timestamp 1751266522
transform 1 0 3516 0 -1 1105
box -2 -3 18 103
use AOI22X1  AOI22X1_44
timestamp 1751266522
transform 1 0 3532 0 -1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_117
timestamp 1751266522
transform -1 0 3604 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_186
timestamp 1751266522
transform -1 0 3628 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_139
timestamp 1751266522
transform 1 0 3628 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_163
timestamp 1751266522
transform -1 0 3668 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_162
timestamp 1751266522
transform -1 0 3692 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_140
timestamp 1751266522
transform -1 0 3708 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_178
timestamp 1751266522
transform -1 0 3732 0 -1 1105
box -2 -3 26 103
use INVX2  INVX2_108
timestamp 1751266522
transform -1 0 3748 0 -1 1105
box -2 -3 18 103
use DFFSR  DFFSR_194
timestamp 1751266522
transform -1 0 3924 0 -1 1105
box -2 -3 178 103
use NAND3X1  NAND3X1_245
timestamp 1751266522
transform 1 0 3924 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_97
timestamp 1751266522
transform -1 0 3988 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_7_0
timestamp 1751266522
transform 1 0 3988 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_7_1
timestamp 1751266522
transform 1 0 3996 0 -1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_95
timestamp 1751266522
transform 1 0 4004 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_102
timestamp 1751266522
transform 1 0 4036 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_168
timestamp 1751266522
transform 1 0 4068 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_33
timestamp 1751266522
transform 1 0 4100 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_247
timestamp 1751266522
transform -1 0 4164 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1751266522
transform 1 0 4164 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_250
timestamp 1751266522
transform 1 0 4196 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_123
timestamp 1751266522
transform 1 0 4228 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1751266522
transform -1 0 4292 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_64
timestamp 1751266522
transform -1 0 4324 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_74
timestamp 1751266522
transform 1 0 4324 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_59
timestamp 1751266522
transform 1 0 4356 0 -1 1105
box -2 -3 34 103
use FILL  FILL_11_1
timestamp 1751266522
transform -1 0 4396 0 -1 1105
box -2 -3 10 103
use BUFX2  BUFX2_82
timestamp 1751266522
transform -1 0 28 0 1 1105
box -2 -3 26 103
use INVX8  INVX8_3
timestamp 1751266522
transform 1 0 28 0 1 1105
box -2 -3 42 103
use BUFX2  BUFX2_7
timestamp 1751266522
transform -1 0 92 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_31
timestamp 1751266522
transform 1 0 92 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_130
timestamp 1751266522
transform 1 0 124 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_209
timestamp 1751266522
transform -1 0 188 0 1 1105
box -2 -3 34 103
use DFFSR  DFFSR_51
timestamp 1751266522
transform 1 0 188 0 1 1105
box -2 -3 178 103
use INVX2  INVX2_3
timestamp 1751266522
transform 1 0 364 0 1 1105
box -2 -3 18 103
use INVX2  INVX2_8
timestamp 1751266522
transform 1 0 380 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_0_0
timestamp 1751266522
transform 1 0 396 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1751266522
transform 1 0 404 0 1 1105
box -2 -3 10 103
use INVX2  INVX2_5
timestamp 1751266522
transform 1 0 412 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_36
timestamp 1751266522
transform -1 0 460 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1751266522
transform 1 0 460 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_40
timestamp 1751266522
transform 1 0 492 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1751266522
transform 1 0 524 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_43
timestamp 1751266522
transform 1 0 556 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_64
timestamp 1751266522
transform 1 0 572 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_100
timestamp 1751266522
transform -1 0 636 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1751266522
transform 1 0 636 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_53
timestamp 1751266522
transform 1 0 668 0 1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_14
timestamp 1751266522
transform -1 0 740 0 1 1105
box -2 -3 42 103
use OAI22X1  OAI22X1_8
timestamp 1751266522
transform 1 0 740 0 1 1105
box -2 -3 42 103
use BUFX4  BUFX4_114
timestamp 1751266522
transform -1 0 812 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_601
timestamp 1751266522
transform 1 0 812 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_59
timestamp 1751266522
transform 1 0 844 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_61
timestamp 1751266522
transform -1 0 892 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1751266522
transform 1 0 892 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1751266522
transform 1 0 900 0 1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_82
timestamp 1751266522
transform 1 0 908 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_61
timestamp 1751266522
transform -1 0 956 0 1 1105
box -2 -3 18 103
use OAI22X1  OAI22X1_43
timestamp 1751266522
transform 1 0 956 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_60
timestamp 1751266522
transform -1 0 1012 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_11
timestamp 1751266522
transform -1 0 1044 0 1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_9
timestamp 1751266522
transform 1 0 1044 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_249
timestamp 1751266522
transform 1 0 1084 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_15
timestamp 1751266522
transform -1 0 1148 0 1 1105
box -2 -3 42 103
use DFFSR  DFFSR_158
timestamp 1751266522
transform 1 0 1148 0 1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_595
timestamp 1751266522
transform 1 0 1324 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1751266522
transform -1 0 1372 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_169
timestamp 1751266522
transform -1 0 1404 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_2_0
timestamp 1751266522
transform 1 0 1404 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1751266522
transform 1 0 1412 0 1 1105
box -2 -3 10 103
use BUFX4  BUFX4_170
timestamp 1751266522
transform 1 0 1420 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_31
timestamp 1751266522
transform 1 0 1452 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_114
timestamp 1751266522
transform 1 0 1492 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_80
timestamp 1751266522
transform -1 0 1540 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_270
timestamp 1751266522
transform 1 0 1540 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_78
timestamp 1751266522
transform 1 0 1572 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_339
timestamp 1751266522
transform 1 0 1604 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_316
timestamp 1751266522
transform 1 0 1636 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_89
timestamp 1751266522
transform 1 0 1668 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_308
timestamp 1751266522
transform 1 0 1692 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_130
timestamp 1751266522
transform 1 0 1724 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_149
timestamp 1751266522
transform 1 0 1740 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_223
timestamp 1751266522
transform 1 0 1756 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_274
timestamp 1751266522
transform -1 0 1820 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_314
timestamp 1751266522
transform 1 0 1820 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_71
timestamp 1751266522
transform -1 0 1876 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_186
timestamp 1751266522
transform -1 0 1900 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_229
timestamp 1751266522
transform -1 0 1924 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_3_0
timestamp 1751266522
transform 1 0 1924 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1751266522
transform 1 0 1932 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_224
timestamp 1751266522
transform 1 0 1940 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_614
timestamp 1751266522
transform 1 0 1964 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_115
timestamp 1751266522
transform 1 0 1996 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_238
timestamp 1751266522
transform -1 0 2188 0 1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_226
timestamp 1751266522
transform -1 0 2212 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_548
timestamp 1751266522
transform 1 0 2212 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_567
timestamp 1751266522
transform 1 0 2244 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_183
timestamp 1751266522
transform 1 0 2276 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_192
timestamp 1751266522
transform 1 0 2308 0 1 1105
box -2 -3 34 103
use DFFSR  DFFSR_186
timestamp 1751266522
transform -1 0 2516 0 1 1105
box -2 -3 178 103
use FILL  FILL_11_4_0
timestamp 1751266522
transform 1 0 2516 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1751266522
transform 1 0 2524 0 1 1105
box -2 -3 10 103
use INVX2  INVX2_114
timestamp 1751266522
transform 1 0 2532 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_691
timestamp 1751266522
transform 1 0 2548 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_219
timestamp 1751266522
transform 1 0 2580 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_78
timestamp 1751266522
transform 1 0 2612 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_187
timestamp 1751266522
transform -1 0 2804 0 1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_171
timestamp 1751266522
transform -1 0 2828 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_97
timestamp 1751266522
transform 1 0 2828 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_488
timestamp 1751266522
transform -1 0 2900 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_487
timestamp 1751266522
transform -1 0 2932 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_486
timestamp 1751266522
transform -1 0 2964 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_5_0
timestamp 1751266522
transform 1 0 2964 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1751266522
transform 1 0 2972 0 1 1105
box -2 -3 10 103
use OAI22X1  OAI22X1_120
timestamp 1751266522
transform 1 0 2980 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_682
timestamp 1751266522
transform -1 0 3052 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_681
timestamp 1751266522
transform -1 0 3084 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_359
timestamp 1751266522
transform -1 0 3116 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_182
timestamp 1751266522
transform 1 0 3116 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_213
timestamp 1751266522
transform 1 0 3140 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_680
timestamp 1751266522
transform -1 0 3204 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_68
timestamp 1751266522
transform 1 0 3204 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_89
timestamp 1751266522
transform 1 0 3220 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_40
timestamp 1751266522
transform 1 0 3252 0 1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_79
timestamp 1751266522
transform 1 0 3292 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_35
timestamp 1751266522
transform 1 0 3324 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_358
timestamp 1751266522
transform 1 0 3364 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_88
timestamp 1751266522
transform -1 0 3428 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_246
timestamp 1751266522
transform -1 0 3460 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_6_0
timestamp 1751266522
transform -1 0 3468 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1751266522
transform -1 0 3476 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_156
timestamp 1751266522
transform -1 0 3500 0 1 1105
box -2 -3 26 103
use INVX2  INVX2_118
timestamp 1751266522
transform 1 0 3500 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_233
timestamp 1751266522
transform -1 0 3692 0 1 1105
box -2 -3 178 103
use INVX1  INVX1_142
timestamp 1751266522
transform -1 0 3708 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_466
timestamp 1751266522
transform -1 0 3740 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_143
timestamp 1751266522
transform 1 0 3740 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_116
timestamp 1751266522
transform -1 0 3788 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_106
timestamp 1751266522
transform 1 0 3788 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_379
timestamp 1751266522
transform -1 0 3836 0 1 1105
box -2 -3 34 103
use AND2X2  AND2X2_15
timestamp 1751266522
transform 1 0 3836 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_109
timestamp 1751266522
transform -1 0 3900 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_108
timestamp 1751266522
transform -1 0 3932 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_141
timestamp 1751266522
transform -1 0 3948 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_99
timestamp 1751266522
transform 1 0 3948 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_7_0
timestamp 1751266522
transform 1 0 3980 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_7_1
timestamp 1751266522
transform 1 0 3988 0 1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_186
timestamp 1751266522
transform 1 0 3996 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_167
timestamp 1751266522
transform 1 0 4028 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_34
timestamp 1751266522
transform 1 0 4060 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_169
timestamp 1751266522
transform -1 0 4124 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_216
timestamp 1751266522
transform 1 0 4124 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_171
timestamp 1751266522
transform 1 0 4156 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_183
timestamp 1751266522
transform 1 0 4188 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_180
timestamp 1751266522
transform 1 0 4220 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_184
timestamp 1751266522
transform -1 0 4284 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_125
timestamp 1751266522
transform 1 0 4284 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_124
timestamp 1751266522
transform 1 0 4316 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_120
timestamp 1751266522
transform 1 0 4348 0 1 1105
box -2 -3 34 103
use FILL  FILL_12_1
timestamp 1751266522
transform 1 0 4380 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1751266522
transform 1 0 4388 0 1 1105
box -2 -3 10 103
use DFFSR  DFFSR_46
timestamp 1751266522
transform -1 0 180 0 -1 1305
box -2 -3 178 103
use DFFSR  DFFSR_61
timestamp 1751266522
transform 1 0 180 0 -1 1305
box -2 -3 178 103
use INVX2  INVX2_37
timestamp 1751266522
transform 1 0 356 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_106
timestamp 1751266522
transform 1 0 372 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1751266522
transform -1 0 412 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1751266522
transform -1 0 420 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_199
timestamp 1751266522
transform -1 0 452 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1751266522
transform 1 0 452 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1751266522
transform 1 0 484 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_22
timestamp 1751266522
transform 1 0 516 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1751266522
transform 1 0 548 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1751266522
transform 1 0 580 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1751266522
transform -1 0 644 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1751266522
transform -1 0 668 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1751266522
transform -1 0 692 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_32
timestamp 1751266522
transform -1 0 716 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_6
timestamp 1751266522
transform -1 0 740 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_41
timestamp 1751266522
transform 1 0 740 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_8
timestamp 1751266522
transform -1 0 788 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_27
timestamp 1751266522
transform -1 0 836 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_49
timestamp 1751266522
transform -1 0 860 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1751266522
transform 1 0 860 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1751266522
transform 1 0 892 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1751266522
transform 1 0 900 0 -1 1305
box -2 -3 10 103
use OAI22X1  OAI22X1_44
timestamp 1751266522
transform 1 0 908 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_31
timestamp 1751266522
transform 1 0 948 0 -1 1305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_31
timestamp 1751266522
transform 1 0 972 0 -1 1305
box -2 -3 74 103
use BUFX4  BUFX4_135
timestamp 1751266522
transform 1 0 1044 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1751266522
transform -1 0 1100 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_192
timestamp 1751266522
transform 1 0 1100 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_85
timestamp 1751266522
transform 1 0 1124 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1751266522
transform 1 0 1156 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_22
timestamp 1751266522
transform -1 0 1220 0 -1 1305
box -2 -3 42 103
use BUFX4  BUFX4_178
timestamp 1751266522
transform -1 0 1252 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_227
timestamp 1751266522
transform -1 0 1284 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1751266522
transform 1 0 1284 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_684
timestamp 1751266522
transform 1 0 1316 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_96
timestamp 1751266522
transform 1 0 1348 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_310
timestamp 1751266522
transform 1 0 1364 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_305
timestamp 1751266522
transform 1 0 1396 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_2_0
timestamp 1751266522
transform 1 0 1428 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1751266522
transform 1 0 1436 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_115
timestamp 1751266522
transform 1 0 1444 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_68
timestamp 1751266522
transform -1 0 1508 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_306
timestamp 1751266522
transform -1 0 1540 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_307
timestamp 1751266522
transform 1 0 1540 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_335
timestamp 1751266522
transform 1 0 1572 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_141
timestamp 1751266522
transform 1 0 1604 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_81
timestamp 1751266522
transform 1 0 1628 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_140
timestamp 1751266522
transform -1 0 1692 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_21
timestamp 1751266522
transform 1 0 1692 0 -1 1305
box -2 -3 42 103
use BUFX4  BUFX4_36
timestamp 1751266522
transform -1 0 1764 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1751266522
transform -1 0 1780 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_46
timestamp 1751266522
transform -1 0 1828 0 -1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_24
timestamp 1751266522
transform -1 0 1876 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_218
timestamp 1751266522
transform 1 0 1876 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_654
timestamp 1751266522
transform 1 0 1900 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1751266522
transform -1 0 1940 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1751266522
transform -1 0 1948 0 -1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_40
timestamp 1751266522
transform -1 0 1996 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_240
timestamp 1751266522
transform -1 0 2020 0 -1 1305
box -2 -3 26 103
use INVX8  INVX8_25
timestamp 1751266522
transform -1 0 2060 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_95
timestamp 1751266522
transform 1 0 2060 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_243
timestamp 1751266522
transform 1 0 2076 0 -1 1305
box -2 -3 26 103
use DFFSR  DFFSR_236
timestamp 1751266522
transform -1 0 2276 0 -1 1305
box -2 -3 178 103
use INVX2  INVX2_139
timestamp 1751266522
transform 1 0 2276 0 -1 1305
box -2 -3 18 103
use INVX4  INVX4_11
timestamp 1751266522
transform 1 0 2292 0 -1 1305
box -2 -3 26 103
use DFFSR  DFFSR_179
timestamp 1751266522
transform -1 0 2492 0 -1 1305
box -2 -3 178 103
use FILL  FILL_12_4_0
timestamp 1751266522
transform 1 0 2492 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1751266522
transform 1 0 2500 0 -1 1305
box -2 -3 10 103
use INVX2  INVX2_116
timestamp 1751266522
transform 1 0 2508 0 -1 1305
box -2 -3 18 103
use DFFSR  DFFSR_174
timestamp 1751266522
transform -1 0 2700 0 -1 1305
box -2 -3 178 103
use AOI22X1  AOI22X1_70
timestamp 1751266522
transform 1 0 2700 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_519
timestamp 1751266522
transform 1 0 2740 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1751266522
transform -1 0 2804 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_67
timestamp 1751266522
transform 1 0 2804 0 -1 1305
box -2 -3 18 103
use DFFSR  DFFSR_211
timestamp 1751266522
transform -1 0 2996 0 -1 1305
box -2 -3 178 103
use FILL  FILL_12_5_0
timestamp 1751266522
transform 1 0 2996 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1751266522
transform 1 0 3004 0 -1 1305
box -2 -3 10 103
use INVX2  INVX2_63
timestamp 1751266522
transform 1 0 3012 0 -1 1305
box -2 -3 18 103
use OAI22X1  OAI22X1_99
timestamp 1751266522
transform 1 0 3028 0 -1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_160
timestamp 1751266522
transform -1 0 3100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_495
timestamp 1751266522
transform 1 0 3100 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_76
timestamp 1751266522
transform 1 0 3132 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_693
timestamp 1751266522
transform -1 0 3180 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1751266522
transform 1 0 3180 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_349
timestamp 1751266522
transform -1 0 3244 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_221
timestamp 1751266522
transform 1 0 3244 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_89
timestamp 1751266522
transform 1 0 3276 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_692
timestamp 1751266522
transform 1 0 3316 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_220
timestamp 1751266522
transform 1 0 3348 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_253
timestamp 1751266522
transform -1 0 3404 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_93
timestamp 1751266522
transform 1 0 3404 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_42
timestamp 1751266522
transform 1 0 3436 0 -1 1305
box -2 -3 42 103
use FILL  FILL_12_6_0
timestamp 1751266522
transform 1 0 3476 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1751266522
transform 1 0 3484 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_346
timestamp 1751266522
transform 1 0 3492 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_78
timestamp 1751266522
transform 1 0 3524 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_265
timestamp 1751266522
transform -1 0 3588 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_16
timestamp 1751266522
transform -1 0 3620 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_156
timestamp 1751266522
transform -1 0 3644 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_245
timestamp 1751266522
transform 1 0 3644 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_155
timestamp 1751266522
transform -1 0 3692 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_366
timestamp 1751266522
transform 1 0 3692 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_96
timestamp 1751266522
transform -1 0 3756 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_157
timestamp 1751266522
transform -1 0 3780 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_362
timestamp 1751266522
transform 1 0 3780 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_92
timestamp 1751266522
transform -1 0 3844 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_268
timestamp 1751266522
transform 1 0 3844 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_160
timestamp 1751266522
transform 1 0 3876 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_106
timestamp 1751266522
transform 1 0 3900 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_107
timestamp 1751266522
transform 1 0 3932 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_7_0
timestamp 1751266522
transform -1 0 3972 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_7_1
timestamp 1751266522
transform -1 0 3980 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_100
timestamp 1751266522
transform -1 0 4012 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_98
timestamp 1751266522
transform 1 0 4012 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_105
timestamp 1751266522
transform 1 0 4044 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_35
timestamp 1751266522
transform 1 0 4076 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_65
timestamp 1751266522
transform 1 0 4108 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_172
timestamp 1751266522
transform 1 0 4140 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_45
timestamp 1751266522
transform 1 0 4172 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_179
timestamp 1751266522
transform 1 0 4204 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_181
timestamp 1751266522
transform -1 0 4268 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_47
timestamp 1751266522
transform 1 0 4268 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1751266522
transform -1 0 4332 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_122
timestamp 1751266522
transform 1 0 4332 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_137
timestamp 1751266522
transform 1 0 4364 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_11
timestamp 1751266522
transform -1 0 28 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_18
timestamp 1751266522
transform -1 0 52 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_141
timestamp 1751266522
transform 1 0 52 0 1 1305
box -2 -3 34 103
use BUFX2  BUFX2_50
timestamp 1751266522
transform -1 0 108 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1751266522
transform 1 0 108 0 1 1305
box -2 -3 34 103
use DFFSR  DFFSR_79
timestamp 1751266522
transform -1 0 316 0 1 1305
box -2 -3 178 103
use FILL  FILL_13_0_0
timestamp 1751266522
transform -1 0 324 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1751266522
transform -1 0 332 0 1 1305
box -2 -3 10 103
use DFFSR  DFFSR_9
timestamp 1751266522
transform -1 0 508 0 1 1305
box -2 -3 178 103
use DFFSR  DFFSR_16
timestamp 1751266522
transform 1 0 508 0 1 1305
box -2 -3 178 103
use NAND2X1  NAND2X1_23
timestamp 1751266522
transform -1 0 708 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1751266522
transform 1 0 708 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_48
timestamp 1751266522
transform 1 0 724 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1751266522
transform 1 0 756 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1751266522
transform 1 0 788 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_47
timestamp 1751266522
transform -1 0 852 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_62
timestamp 1751266522
transform 1 0 852 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_113
timestamp 1751266522
transform 1 0 884 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1751266522
transform 1 0 916 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1751266522
transform 1 0 924 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_39
timestamp 1751266522
transform 1 0 932 0 1 1305
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1751266522
transform 1 0 964 0 1 1305
box -2 -3 42 103
use BUFX4  BUFX4_192
timestamp 1751266522
transform 1 0 1004 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_24
timestamp 1751266522
transform 1 0 1036 0 1 1305
box -2 -3 42 103
use INVX1  INVX1_41
timestamp 1751266522
transform -1 0 1092 0 1 1305
box -2 -3 18 103
use OAI22X1  OAI22X1_21
timestamp 1751266522
transform -1 0 1132 0 1 1305
box -2 -3 42 103
use INVX1  INVX1_38
timestamp 1751266522
transform -1 0 1148 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_31
timestamp 1751266522
transform 1 0 1148 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_629
timestamp 1751266522
transform 1 0 1196 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_46
timestamp 1751266522
transform 1 0 1228 0 1 1305
box -2 -3 42 103
use BUFX4  BUFX4_239
timestamp 1751266522
transform -1 0 1300 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_177
timestamp 1751266522
transform 1 0 1300 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_49
timestamp 1751266522
transform -1 0 1340 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_19
timestamp 1751266522
transform 1 0 1340 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_586
timestamp 1751266522
transform 1 0 1388 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_2_0
timestamp 1751266522
transform -1 0 1428 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1751266522
transform -1 0 1436 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_63
timestamp 1751266522
transform -1 0 1452 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_628
timestamp 1751266522
transform 1 0 1452 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_242
timestamp 1751266522
transform 1 0 1484 0 1 1305
box -2 -3 34 103
use INVX8  INVX8_6
timestamp 1751266522
transform 1 0 1516 0 1 1305
box -2 -3 42 103
use INVX1  INVX1_50
timestamp 1751266522
transform -1 0 1572 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_119
timestamp 1751266522
transform 1 0 1572 0 1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_70
timestamp 1751266522
transform -1 0 1636 0 1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_118
timestamp 1751266522
transform 1 0 1636 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_311
timestamp 1751266522
transform -1 0 1692 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_142
timestamp 1751266522
transform 1 0 1692 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_312
timestamp 1751266522
transform -1 0 1748 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_69
timestamp 1751266522
transform 1 0 1748 0 1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_116
timestamp 1751266522
transform -1 0 1812 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_341
timestamp 1751266522
transform 1 0 1812 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_112
timestamp 1751266522
transform 1 0 1844 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_340
timestamp 1751266522
transform -1 0 1892 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_300
timestamp 1751266522
transform 1 0 1892 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_3_0
timestamp 1751266522
transform -1 0 1932 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1751266522
transform -1 0 1940 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_34
timestamp 1751266522
transform -1 0 1972 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_109
timestamp 1751266522
transform 1 0 1972 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_249
timestamp 1751266522
transform 1 0 1988 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_32
timestamp 1751266522
transform -1 0 2060 0 1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_251
timestamp 1751266522
transform -1 0 2084 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_234
timestamp 1751266522
transform 1 0 2084 0 1 1305
box -2 -3 26 103
use DFFSR  DFFSR_119
timestamp 1751266522
transform -1 0 2284 0 1 1305
box -2 -3 178 103
use OAI21X1  OAI21X1_594
timestamp 1751266522
transform 1 0 2284 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_683
timestamp 1751266522
transform 1 0 2316 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_119
timestamp 1751266522
transform 1 0 2348 0 1 1305
box -2 -3 18 103
use AOI22X1  AOI22X1_75
timestamp 1751266522
transform 1 0 2364 0 1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_188
timestamp 1751266522
transform -1 0 2436 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_4_0
timestamp 1751266522
transform -1 0 2444 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1751266522
transform -1 0 2452 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_559
timestamp 1751266522
transform -1 0 2484 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_69
timestamp 1751266522
transform 1 0 2484 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_187
timestamp 1751266522
transform 1 0 2500 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_558
timestamp 1751266522
transform -1 0 2564 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_672
timestamp 1751266522
transform 1 0 2564 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_210
timestamp 1751266522
transform 1 0 2596 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_84
timestamp 1751266522
transform 1 0 2628 0 1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_671
timestamp 1751266522
transform 1 0 2668 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_209
timestamp 1751266522
transform -1 0 2732 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_248
timestamp 1751266522
transform -1 0 2756 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_169
timestamp 1751266522
transform -1 0 2788 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_212
timestamp 1751266522
transform -1 0 2812 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_520
timestamp 1751266522
transform -1 0 2844 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_664
timestamp 1751266522
transform -1 0 2876 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_204
timestamp 1751266522
transform 1 0 2876 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_118
timestamp 1751266522
transform -1 0 2948 0 1 1305
box -2 -3 42 103
use FILL  FILL_13_5_0
timestamp 1751266522
transform -1 0 2956 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1751266522
transform -1 0 2964 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_666
timestamp 1751266522
transform -1 0 2996 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_665
timestamp 1751266522
transform -1 0 3028 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1751266522
transform -1 0 3060 0 1 1305
box -2 -3 34 103
use DFFSR  DFFSR_219
timestamp 1751266522
transform -1 0 3236 0 1 1305
box -2 -3 178 103
use OAI21X1  OAI21X1_363
timestamp 1751266522
transform -1 0 3268 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_154
timestamp 1751266522
transform -1 0 3284 0 1 1305
box -2 -3 18 103
use BUFX4  BUFX4_253
timestamp 1751266522
transform -1 0 3316 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_396
timestamp 1751266522
transform -1 0 3348 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_112
timestamp 1751266522
transform -1 0 3364 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_388
timestamp 1751266522
transform -1 0 3396 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_184
timestamp 1751266522
transform -1 0 3420 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_6_0
timestamp 1751266522
transform -1 0 3428 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1751266522
transform -1 0 3436 0 1 1305
box -2 -3 10 103
use DFFSR  DFFSR_218
timestamp 1751266522
transform -1 0 3612 0 1 1305
box -2 -3 178 103
use NAND2X1  NAND2X1_133
timestamp 1751266522
transform -1 0 3636 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_123
timestamp 1751266522
transform 1 0 3636 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_54
timestamp 1751266522
transform 1 0 3668 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_164
timestamp 1751266522
transform 1 0 3708 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_160
timestamp 1751266522
transform 1 0 3732 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_153
timestamp 1751266522
transform -1 0 3772 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_160
timestamp 1751266522
transform 1 0 3772 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_191
timestamp 1751266522
transform -1 0 3820 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_395
timestamp 1751266522
transform 1 0 3820 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_122
timestamp 1751266522
transform -1 0 3884 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_227
timestamp 1751266522
transform 1 0 3884 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_192
timestamp 1751266522
transform 1 0 3916 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_108
timestamp 1751266522
transform 1 0 3948 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_7_0
timestamp 1751266522
transform 1 0 3980 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_7_1
timestamp 1751266522
transform 1 0 3988 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_36
timestamp 1751266522
transform 1 0 3996 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_193
timestamp 1751266522
transform 1 0 4028 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_189
timestamp 1751266522
transform 1 0 4060 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_217
timestamp 1751266522
transform 1 0 4092 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_170
timestamp 1751266522
transform 1 0 4124 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_187
timestamp 1751266522
transform 1 0 4156 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_224
timestamp 1751266522
transform 1 0 4188 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_188
timestamp 1751266522
transform -1 0 4252 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_225
timestamp 1751266522
transform 1 0 4252 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_185
timestamp 1751266522
transform -1 0 4316 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_219
timestamp 1751266522
transform 1 0 4316 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_205
timestamp 1751266522
transform 1 0 4348 0 1 1305
box -2 -3 34 103
use FILL  FILL_14_1
timestamp 1751266522
transform 1 0 4380 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1751266522
transform 1 0 4388 0 1 1305
box -2 -3 10 103
use BUFX2  BUFX2_10
timestamp 1751266522
transform -1 0 28 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_133
timestamp 1751266522
transform -1 0 60 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_17
timestamp 1751266522
transform 1 0 60 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_8
timestamp 1751266522
transform -1 0 252 0 -1 1505
box -2 -3 178 103
use BUFX4  BUFX4_208
timestamp 1751266522
transform 1 0 252 0 -1 1505
box -2 -3 34 103
use DFFSR  DFFSR_49
timestamp 1751266522
transform 1 0 284 0 -1 1505
box -2 -3 178 103
use FILL  FILL_14_0_0
timestamp 1751266522
transform 1 0 460 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1751266522
transform 1 0 468 0 -1 1505
box -2 -3 10 103
use INVX2  INVX2_2
timestamp 1751266522
transform 1 0 476 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_64
timestamp 1751266522
transform -1 0 524 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1751266522
transform 1 0 524 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1751266522
transform 1 0 556 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1751266522
transform 1 0 588 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_101
timestamp 1751266522
transform -1 0 652 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_63
timestamp 1751266522
transform 1 0 652 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_103
timestamp 1751266522
transform 1 0 684 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_23
timestamp 1751266522
transform 1 0 716 0 -1 1505
box -2 -3 42 103
use BUFX4  BUFX4_96
timestamp 1751266522
transform -1 0 788 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_194
timestamp 1751266522
transform -1 0 820 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1751266522
transform -1 0 844 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_245
timestamp 1751266522
transform -1 0 868 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_1
timestamp 1751266522
transform 1 0 868 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_1_0
timestamp 1751266522
transform -1 0 908 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1751266522
transform -1 0 916 0 -1 1505
box -2 -3 10 103
use INVX2  INVX2_1
timestamp 1751266522
transform -1 0 932 0 -1 1505
box -2 -3 18 103
use BUFX4  BUFX4_133
timestamp 1751266522
transform -1 0 964 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_69
timestamp 1751266522
transform -1 0 996 0 -1 1505
box -2 -3 34 103
use INVX4  INVX4_1
timestamp 1751266522
transform -1 0 1020 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_71
timestamp 1751266522
transform -1 0 1052 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1751266522
transform -1 0 1076 0 -1 1505
box -2 -3 26 103
use DFFSR  DFFSR_130
timestamp 1751266522
transform -1 0 1252 0 -1 1505
box -2 -3 178 103
use AOI21X1  AOI21X1_18
timestamp 1751266522
transform -1 0 1284 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1751266522
transform 1 0 1284 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_31
timestamp 1751266522
transform 1 0 1316 0 -1 1505
box -2 -3 42 103
use OAI22X1  OAI22X1_10
timestamp 1751266522
transform -1 0 1396 0 -1 1505
box -2 -3 42 103
use INVX1  INVX1_27
timestamp 1751266522
transform -1 0 1412 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_2_0
timestamp 1751266522
transform -1 0 1420 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1751266522
transform -1 0 1428 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_151
timestamp 1751266522
transform -1 0 1452 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_25
timestamp 1751266522
transform -1 0 1476 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_48
timestamp 1751266522
transform -1 0 1492 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_28
timestamp 1751266522
transform 1 0 1492 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_20
timestamp 1751266522
transform -1 0 1540 0 -1 1505
box -2 -3 26 103
use INVX8  INVX8_15
timestamp 1751266522
transform 1 0 1540 0 -1 1505
box -2 -3 42 103
use OAI22X1  OAI22X1_52
timestamp 1751266522
transform -1 0 1620 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_79
timestamp 1751266522
transform 1 0 1620 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_263
timestamp 1751266522
transform -1 0 1676 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_51
timestamp 1751266522
transform -1 0 1716 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_77
timestamp 1751266522
transform 1 0 1716 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_117
timestamp 1751266522
transform -1 0 1764 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_87
timestamp 1751266522
transform 1 0 1764 0 -1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_55
timestamp 1751266522
transform -1 0 1828 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_86
timestamp 1751266522
transform -1 0 1852 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_142
timestamp 1751266522
transform -1 0 1876 0 -1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_82
timestamp 1751266522
transform 1 0 1876 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_143
timestamp 1751266522
transform -1 0 1940 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_3_0
timestamp 1751266522
transform 1 0 1940 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1751266522
transform 1 0 1948 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_39
timestamp 1751266522
transform 1 0 1956 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_655
timestamp 1751266522
transform -1 0 2036 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_275
timestamp 1751266522
transform 1 0 2036 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_255
timestamp 1751266522
transform 1 0 2068 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_695
timestamp 1751266522
transform -1 0 2124 0 -1 1505
box -2 -3 34 103
use DFFSR  DFFSR_131
timestamp 1751266522
transform -1 0 2300 0 -1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_696
timestamp 1751266522
transform 1 0 2300 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1751266522
transform -1 0 2364 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1751266522
transform -1 0 2396 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_219
timestamp 1751266522
transform 1 0 2396 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_217
timestamp 1751266522
transform 1 0 2420 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_4_0
timestamp 1751266522
transform 1 0 2444 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1751266522
transform 1 0 2452 0 -1 1505
box -2 -3 10 103
use INVX2  INVX2_71
timestamp 1751266522
transform 1 0 2460 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_163
timestamp 1751266522
transform -1 0 2652 0 -1 1505
box -2 -3 178 103
use AOI22X1  AOI22X1_86
timestamp 1751266522
transform 1 0 2652 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_250
timestamp 1751266522
transform 1 0 2692 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_686
timestamp 1751266522
transform 1 0 2716 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_214
timestamp 1751266522
transform 1 0 2748 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_201
timestamp 1751266522
transform 1 0 2780 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_195
timestamp 1751266522
transform 1 0 2804 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_246
timestamp 1751266522
transform 1 0 2828 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_244
timestamp 1751266522
transform 1 0 2852 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_5_0
timestamp 1751266522
transform -1 0 2884 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1751266522
transform -1 0 2892 0 -1 1505
box -2 -3 10 103
use DFFSR  DFFSR_183
timestamp 1751266522
transform -1 0 3068 0 -1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_427
timestamp 1751266522
transform -1 0 3100 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_117
timestamp 1751266522
transform -1 0 3116 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_206
timestamp 1751266522
transform -1 0 3292 0 -1 1505
box -2 -3 178 103
use NOR2X1  NOR2X1_177
timestamp 1751266522
transform -1 0 3316 0 -1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_86
timestamp 1751266522
transform 1 0 3316 0 -1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_428
timestamp 1751266522
transform -1 0 3388 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_140
timestamp 1751266522
transform -1 0 3420 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_426
timestamp 1751266522
transform -1 0 3452 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_168
timestamp 1751266522
transform 1 0 3452 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_6_0
timestamp 1751266522
transform -1 0 3484 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1751266522
transform -1 0 3492 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_425
timestamp 1751266522
transform -1 0 3524 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_55
timestamp 1751266522
transform -1 0 3556 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_441
timestamp 1751266522
transform 1 0 3556 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_145
timestamp 1751266522
transform 1 0 3588 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_663
timestamp 1751266522
transform 1 0 3612 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_52
timestamp 1751266522
transform -1 0 3676 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_244
timestamp 1751266522
transform -1 0 3700 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_75
timestamp 1751266522
transform 1 0 3700 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_154
timestamp 1751266522
transform -1 0 3748 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_146
timestamp 1751266522
transform -1 0 3772 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_159
timestamp 1751266522
transform 1 0 3772 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_160
timestamp 1751266522
transform 1 0 3796 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_201
timestamp 1751266522
transform 1 0 3828 0 -1 1505
box -2 -3 26 103
use DFFSR  DFFSR_195
timestamp 1751266522
transform -1 0 4028 0 -1 1505
box -2 -3 178 103
use FILL  FILL_14_7_0
timestamp 1751266522
transform -1 0 4036 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_7_1
timestamp 1751266522
transform -1 0 4044 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_194
timestamp 1751266522
transform -1 0 4076 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_195
timestamp 1751266522
transform 1 0 4076 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_197
timestamp 1751266522
transform 1 0 4108 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_49
timestamp 1751266522
transform 1 0 4140 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_191
timestamp 1751266522
transform 1 0 4172 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_190
timestamp 1751266522
transform 1 0 4204 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1751266522
transform 1 0 4236 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_226
timestamp 1751266522
transform 1 0 4268 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_76
timestamp 1751266522
transform -1 0 4332 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1751266522
transform -1 0 4364 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1751266522
transform -1 0 4396 0 -1 1505
box -2 -3 34 103
use BUFX2  BUFX2_16
timestamp 1751266522
transform -1 0 28 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_32
timestamp 1751266522
transform -1 0 52 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_155
timestamp 1751266522
transform 1 0 52 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_27
timestamp 1751266522
transform 1 0 84 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_139
timestamp 1751266522
transform 1 0 116 0 1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_58
timestamp 1751266522
transform 1 0 148 0 1 1505
box -2 -3 74 103
use BUFX2  BUFX2_30
timestamp 1751266522
transform -1 0 28 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_46
timestamp 1751266522
transform -1 0 52 0 -1 1705
box -2 -3 26 103
use DFFSR  DFFSR_75
timestamp 1751266522
transform -1 0 228 0 -1 1705
box -2 -3 178 103
use DFFSR  DFFSR_14
timestamp 1751266522
transform -1 0 396 0 1 1505
box -2 -3 178 103
use BUFX4  BUFX4_215
timestamp 1751266522
transform 1 0 228 0 -1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1751266522
transform -1 0 332 0 -1 1705
box -2 -3 74 103
use BUFX4  BUFX4_29
timestamp 1751266522
transform -1 0 364 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1751266522
transform 1 0 364 0 -1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_23
timestamp 1751266522
transform 1 0 412 0 -1 1705
box -2 -3 74 103
use FILL  FILL_16_0_1
timestamp 1751266522
transform 1 0 404 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_0
timestamp 1751266522
transform 1 0 396 0 -1 1705
box -2 -3 10 103
use BUFX4  BUFX4_118
timestamp 1751266522
transform -1 0 460 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_7
timestamp 1751266522
transform 1 0 412 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_0_1
timestamp 1751266522
transform 1 0 404 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_0
timestamp 1751266522
transform 1 0 396 0 1 1505
box -2 -3 10 103
use INVX2  INVX2_16
timestamp 1751266522
transform 1 0 484 0 -1 1705
box -2 -3 18 103
use DFFSR  DFFSR_28
timestamp 1751266522
transform -1 0 676 0 -1 1705
box -2 -3 178 103
use DFFSR  DFFSR_56
timestamp 1751266522
transform 1 0 460 0 1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_44
timestamp 1751266522
transform 1 0 636 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_32
timestamp 1751266522
transform 1 0 668 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_96
timestamp 1751266522
transform 1 0 684 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_201
timestamp 1751266522
transform -1 0 748 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_62
timestamp 1751266522
transform 1 0 676 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1751266522
transform 1 0 708 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1751266522
transform 1 0 772 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1751266522
transform 1 0 740 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_53
timestamp 1751266522
transform 1 0 748 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1751266522
transform 1 0 804 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1751266522
transform -1 0 844 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1751266522
transform 1 0 780 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_50
timestamp 1751266522
transform 1 0 836 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_33
timestamp 1751266522
transform -1 0 876 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1_0
timestamp 1751266522
transform -1 0 908 0 -1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_27
timestamp 1751266522
transform -1 0 900 0 -1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_29
timestamp 1751266522
transform -1 0 916 0 1 1505
box -2 -3 42 103
use FILL  FILL_16_1_1
timestamp 1751266522
transform -1 0 916 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_61
timestamp 1751266522
transform 1 0 948 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1751266522
transform -1 0 948 0 -1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_20
timestamp 1751266522
transform 1 0 932 0 1 1505
box -2 -3 42 103
use FILL  FILL_15_1_1
timestamp 1751266522
transform 1 0 924 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_0
timestamp 1751266522
transform 1 0 916 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_97
timestamp 1751266522
transform -1 0 1012 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_217
timestamp 1751266522
transform -1 0 1004 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1751266522
transform 1 0 1012 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_19
timestamp 1751266522
transform 1 0 1036 0 1 1505
box -2 -3 18 103
use BUFX4  BUFX4_219
timestamp 1751266522
transform -1 0 1036 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1751266522
transform -1 0 1100 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1751266522
transform 1 0 1044 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_35
timestamp 1751266522
transform 1 0 1084 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_51
timestamp 1751266522
transform 1 0 1052 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1751266522
transform -1 0 1148 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1751266522
transform 1 0 1100 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_125
timestamp 1751266522
transform 1 0 1116 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_99
timestamp 1751266522
transform 1 0 1148 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_70
timestamp 1751266522
transform 1 0 1148 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1751266522
transform -1 0 1228 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1751266522
transform 1 0 1180 0 -1 1705
box -2 -3 26 103
use INVX8  INVX8_5
timestamp 1751266522
transform 1 0 1212 0 1 1505
box -2 -3 42 103
use NAND3X1  NAND3X1_68
timestamp 1751266522
transform 1 0 1180 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_50
timestamp 1751266522
transform -1 0 1284 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_81
timestamp 1751266522
transform -1 0 1260 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1751266522
transform 1 0 1252 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1751266522
transform 1 0 1308 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1751266522
transform -1 0 1308 0 -1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_33
timestamp 1751266522
transform 1 0 1284 0 1 1505
box -2 -3 42 103
use BUFX4  BUFX4_68
timestamp 1751266522
transform 1 0 1356 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1751266522
transform -1 0 1356 0 -1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_12
timestamp 1751266522
transform -1 0 1396 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_4
timestamp 1751266522
transform 1 0 1324 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_45
timestamp 1751266522
transform 1 0 1388 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_29
timestamp 1751266522
transform -1 0 1412 0 1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_17
timestamp 1751266522
transform -1 0 1476 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_2_1
timestamp 1751266522
transform -1 0 1444 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_0
timestamp 1751266522
transform -1 0 1436 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_585
timestamp 1751266522
transform 1 0 1444 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_62
timestamp 1751266522
transform -1 0 1444 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_2_1
timestamp 1751266522
transform -1 0 1428 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_0
timestamp 1751266522
transform -1 0 1420 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_132
timestamp 1751266522
transform 1 0 1476 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_163
timestamp 1751266522
transform -1 0 1508 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_4
timestamp 1751266522
transform 1 0 1540 0 -1 1705
box -2 -3 42 103
use BUFX4  BUFX4_134
timestamp 1751266522
transform 1 0 1508 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_650
timestamp 1751266522
transform 1 0 1556 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_37
timestamp 1751266522
transform -1 0 1556 0 1 1505
box -2 -3 50 103
use OAI22X1  OAI22X1_25
timestamp 1751266522
transform 1 0 1596 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_22
timestamp 1751266522
transform -1 0 1596 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_649
timestamp 1751266522
transform 1 0 1588 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_21
timestamp 1751266522
transform -1 0 1636 0 1 1505
box -2 -3 18 103
use INVX8  INVX8_7
timestamp 1751266522
transform 1 0 1668 0 -1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_261
timestamp 1751266522
transform -1 0 1668 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_271
timestamp 1751266522
transform 1 0 1668 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_342
timestamp 1751266522
transform -1 0 1668 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_177
timestamp 1751266522
transform 1 0 1708 0 -1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_56
timestamp 1751266522
transform -1 0 1740 0 1 1505
box -2 -3 42 103
use BUFX4  BUFX4_37
timestamp 1751266522
transform -1 0 1796 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_88
timestamp 1751266522
transform 1 0 1740 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_258
timestamp 1751266522
transform 1 0 1740 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_299
timestamp 1751266522
transform -1 0 1828 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_273
timestamp 1751266522
transform 1 0 1804 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_309
timestamp 1751266522
transform -1 0 1804 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1751266522
transform -1 0 1860 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_42
timestamp 1751266522
transform -1 0 1844 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_269
timestamp 1751266522
transform -1 0 1868 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_66
timestamp 1751266522
transform 1 0 1884 0 -1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_109
timestamp 1751266522
transform -1 0 1884 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_343
timestamp 1751266522
transform 1 0 1900 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_171
timestamp 1751266522
transform -1 0 1900 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_226
timestamp 1751266522
transform 1 0 1940 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_3_1
timestamp 1751266522
transform 1 0 1932 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_0
timestamp 1751266522
transform 1 0 1924 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_145
timestamp 1751266522
transform 1 0 1948 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_3_1
timestamp 1751266522
transform 1 0 1940 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_0
timestamp 1751266522
transform 1 0 1932 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_141
timestamp 1751266522
transform 1 0 1972 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_344
timestamp 1751266522
transform 1 0 1972 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1751266522
transform -1 0 2092 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_17
timestamp 1751266522
transform 1 0 2028 0 -1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_301
timestamp 1751266522
transform -1 0 2028 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_238
timestamp 1751266522
transform -1 0 2092 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_38
timestamp 1751266522
transform -1 0 2068 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_106
timestamp 1751266522
transform 1 0 2004 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_323
timestamp 1751266522
transform 1 0 2140 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_146
timestamp 1751266522
transform -1 0 2140 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_194
timestamp 1751266522
transform -1 0 2116 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_640
timestamp 1751266522
transform 1 0 2156 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_639
timestamp 1751266522
transform 1 0 2124 0 1 1505
box -2 -3 34 103
use AND2X2  AND2X2_27
timestamp 1751266522
transform 1 0 2092 0 1 1505
box -2 -3 34 103
use DFFSR  DFFSR_126
timestamp 1751266522
transform -1 0 2348 0 -1 1705
box -2 -3 178 103
use INVX1  INVX1_113
timestamp 1751266522
transform 1 0 2188 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_638
timestamp 1751266522
transform 1 0 2204 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_237
timestamp 1751266522
transform -1 0 2260 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_97
timestamp 1751266522
transform 1 0 2260 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_694
timestamp 1751266522
transform 1 0 2276 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1751266522
transform -1 0 2332 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_153
timestamp 1751266522
transform -1 0 2508 0 1 1505
box -2 -3 178 103
use INVX2  INVX2_101
timestamp 1751266522
transform 1 0 2348 0 -1 1705
box -2 -3 18 103
use FILL  FILL_15_4_0
timestamp 1751266522
transform 1 0 2508 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_1
timestamp 1751266522
transform 1 0 2516 0 1 1505
box -2 -3 10 103
use INVX4  INVX4_12
timestamp 1751266522
transform 1 0 2524 0 1 1505
box -2 -3 26 103
use INVX2  INVX2_95
timestamp 1751266522
transform 1 0 2364 0 -1 1705
box -2 -3 18 103
use FILL  FILL_16_4_0
timestamp 1751266522
transform -1 0 2388 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_1
timestamp 1751266522
transform -1 0 2396 0 -1 1705
box -2 -3 10 103
use DFFSR  DFFSR_149
timestamp 1751266522
transform -1 0 2572 0 -1 1705
box -2 -3 178 103
use INVX1  INVX1_104
timestamp 1751266522
transform 1 0 2572 0 -1 1705
box -2 -3 18 103
use AOI22X1  AOI22X1_77
timestamp 1751266522
transform 1 0 2548 0 1 1505
box -2 -3 42 103
use OAI22X1  OAI22X1_117
timestamp 1751266522
transform 1 0 2588 0 -1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_193
timestamp 1751266522
transform 1 0 2620 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_568
timestamp 1751266522
transform 1 0 2588 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_577
timestamp 1751266522
transform -1 0 2692 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_578
timestamp 1751266522
transform -1 0 2660 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1751266522
transform -1 0 2684 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_569
timestamp 1751266522
transform -1 0 2748 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_212
timestamp 1751266522
transform 1 0 2692 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_687
timestamp 1751266522
transform -1 0 2748 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_215
timestamp 1751266522
transform -1 0 2716 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1751266522
transform 1 0 2748 0 1 1505
box -2 -3 34 103
use DFFSR  DFFSR_181
timestamp 1751266522
transform -1 0 2956 0 1 1505
box -2 -3 178 103
use INVX2  INVX2_72
timestamp 1751266522
transform 1 0 2748 0 -1 1705
box -2 -3 18 103
use BUFX4  BUFX4_150
timestamp 1751266522
transform 1 0 2764 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_526
timestamp 1751266522
transform 1 0 2796 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_525
timestamp 1751266522
transform -1 0 2860 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_140
timestamp 1751266522
transform -1 0 2876 0 -1 1705
box -2 -3 18 103
use CLKBUF1  CLKBUF1_40
timestamp 1751266522
transform -1 0 2948 0 -1 1705
box -2 -3 74 103
use FILL  FILL_15_5_0
timestamp 1751266522
transform 1 0 2956 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_1
timestamp 1751266522
transform 1 0 2964 0 1 1505
box -2 -3 10 103
use DFFSR  DFFSR_213
timestamp 1751266522
transform 1 0 2972 0 1 1505
box -2 -3 178 103
use FILL  FILL_16_5_0
timestamp 1751266522
transform 1 0 2948 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_5_1
timestamp 1751266522
transform 1 0 2956 0 -1 1705
box -2 -3 10 103
use INVX2  INVX2_120
timestamp 1751266522
transform 1 0 2964 0 -1 1705
box -2 -3 18 103
use DFFSR  DFFSR_190
timestamp 1751266522
transform -1 0 3156 0 -1 1705
box -2 -3 178 103
use INVX2  INVX2_96
timestamp 1751266522
transform 1 0 3148 0 1 1505
box -2 -3 18 103
use INVX2  INVX2_94
timestamp 1751266522
transform 1 0 3164 0 1 1505
box -2 -3 18 103
use BUFX4  BUFX4_42
timestamp 1751266522
transform 1 0 3180 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_229
timestamp 1751266522
transform -1 0 3244 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_234
timestamp 1751266522
transform -1 0 3276 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_141
timestamp 1751266522
transform 1 0 3156 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_435
timestamp 1751266522
transform 1 0 3172 0 -1 1705
box -2 -3 34 103
use DFFSR  DFFSR_204
timestamp 1751266522
transform -1 0 3380 0 -1 1705
box -2 -3 178 103
use OAI21X1  OAI21X1_503
timestamp 1751266522
transform 1 0 3276 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_502
timestamp 1751266522
transform -1 0 3340 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_406
timestamp 1751266522
transform -1 0 3372 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_101
timestamp 1751266522
transform 1 0 3372 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_162
timestamp 1751266522
transform 1 0 3412 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_233
timestamp 1751266522
transform 1 0 3380 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_348
timestamp 1751266522
transform 1 0 3412 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_6_1
timestamp 1751266522
transform 1 0 3484 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_0
timestamp 1751266522
transform 1 0 3476 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_668
timestamp 1751266522
transform 1 0 3444 0 -1 1705
box -2 -3 34 103
use FILL  FILL_15_6_1
timestamp 1751266522
transform -1 0 3492 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_6_0
timestamp 1751266522
transform -1 0 3484 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_501
timestamp 1751266522
transform 1 0 3444 0 1 1505
box -2 -3 34 103
use AOI22X1  AOI22X1_82
timestamp 1751266522
transform 1 0 3524 0 -1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_206
timestamp 1751266522
transform 1 0 3492 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_133
timestamp 1751266522
transform 1 0 3516 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_158
timestamp 1751266522
transform -1 0 3516 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_667
timestamp 1751266522
transform 1 0 3564 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_59
timestamp 1751266522
transform 1 0 3548 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_205
timestamp 1751266522
transform -1 0 3628 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_674
timestamp 1751266522
transform -1 0 3644 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_247
timestamp 1751266522
transform 1 0 3588 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_96
timestamp 1751266522
transform -1 0 3740 0 -1 1705
box -2 -3 42 103
use INVX2  INVX2_144
timestamp 1751266522
transform -1 0 3700 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_485
timestamp 1751266522
transform 1 0 3652 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_193
timestamp 1751266522
transform -1 0 3652 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_673
timestamp 1751266522
transform -1 0 3724 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_675
timestamp 1751266522
transform 1 0 3660 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_70
timestamp 1751266522
transform -1 0 3660 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_150
timestamp 1751266522
transform 1 0 3796 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_119
timestamp 1751266522
transform -1 0 3796 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_211
timestamp 1751266522
transform 1 0 3724 0 1 1505
box -2 -3 34 103
use DFFSR  DFFSR_188
timestamp 1751266522
transform -1 0 3916 0 -1 1705
box -2 -3 178 103
use BUFX4  BUFX4_17
timestamp 1751266522
transform 1 0 3820 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_405
timestamp 1751266522
transform 1 0 3852 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_132
timestamp 1751266522
transform -1 0 3916 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_231
timestamp 1751266522
transform 1 0 3948 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_110
timestamp 1751266522
transform 1 0 3916 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_109
timestamp 1751266522
transform 1 0 3932 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_157
timestamp 1751266522
transform -1 0 3932 0 1 1505
box -2 -3 18 103
use FILL  FILL_16_7_0
timestamp 1751266522
transform 1 0 3980 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_37
timestamp 1751266522
transform 1 0 3980 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_7_1
timestamp 1751266522
transform 1 0 3972 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_7_0
timestamp 1751266522
transform 1 0 3964 0 1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_153
timestamp 1751266522
transform 1 0 3996 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_7_1
timestamp 1751266522
transform 1 0 3988 0 -1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_229
timestamp 1751266522
transform 1 0 4012 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_228
timestamp 1751266522
transform 1 0 4028 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_111
timestamp 1751266522
transform 1 0 4044 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_112
timestamp 1751266522
transform 1 0 4092 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_232
timestamp 1751266522
transform -1 0 4092 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1751266522
transform 1 0 4076 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_196
timestamp 1751266522
transform 1 0 4124 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_218
timestamp 1751266522
transform 1 0 4108 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_138
timestamp 1751266522
transform 1 0 4156 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_113
timestamp 1751266522
transform -1 0 4172 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_140
timestamp 1751266522
transform 1 0 4188 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_139
timestamp 1751266522
transform 1 0 4172 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1751266522
transform 1 0 4220 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_137
timestamp 1751266522
transform 1 0 4236 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_135
timestamp 1751266522
transform 1 0 4204 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_136
timestamp 1751266522
transform 1 0 4252 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_142
timestamp 1751266522
transform 1 0 4268 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_141
timestamp 1751266522
transform 1 0 4284 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_210
timestamp 1751266522
transform -1 0 4332 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_59
timestamp 1751266522
transform -1 0 4348 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_126
timestamp 1751266522
transform 1 0 4332 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1
timestamp 1751266522
transform 1 0 4364 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1751266522
transform 1 0 4372 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_3
timestamp 1751266522
transform 1 0 4380 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_4
timestamp 1751266522
transform 1 0 4388 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_229
timestamp 1751266522
transform 1 0 4348 0 -1 1705
box -2 -3 34 103
use FILL  FILL_17_1
timestamp 1751266522
transform -1 0 4388 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_2
timestamp 1751266522
transform -1 0 4396 0 -1 1705
box -2 -3 10 103
use BUFX2  BUFX2_3
timestamp 1751266522
transform -1 0 28 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_65
timestamp 1751266522
transform -1 0 52 0 1 1705
box -2 -3 26 103
use DFFSR  DFFSR_94
timestamp 1751266522
transform -1 0 228 0 1 1705
box -2 -3 178 103
use DFFSR  DFFSR_4
timestamp 1751266522
transform -1 0 404 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_0_0
timestamp 1751266522
transform 1 0 404 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1751266522
transform 1 0 412 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_126
timestamp 1751266522
transform 1 0 420 0 1 1705
box -2 -3 34 103
use DFFSR  DFFSR_7
timestamp 1751266522
transform -1 0 628 0 1 1705
box -2 -3 178 103
use DFFSR  DFFSR_1
timestamp 1751266522
transform 1 0 628 0 1 1705
box -2 -3 178 103
use INVX2  INVX2_10
timestamp 1751266522
transform 1 0 804 0 1 1705
box -2 -3 18 103
use OAI22X1  OAI22X1_11
timestamp 1751266522
transform -1 0 860 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_129
timestamp 1751266522
transform -1 0 892 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_1_0
timestamp 1751266522
transform -1 0 900 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1751266522
transform -1 0 908 0 1 1705
box -2 -3 10 103
use OAI22X1  OAI22X1_26
timestamp 1751266522
transform -1 0 948 0 1 1705
box -2 -3 42 103
use INVX8  INVX8_4
timestamp 1751266522
transform 1 0 948 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_218
timestamp 1751266522
transform -1 0 1020 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_191
timestamp 1751266522
transform -1 0 1052 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1751266522
transform 1 0 1052 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1751266522
transform 1 0 1084 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_193
timestamp 1751266522
transform 1 0 1116 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_198
timestamp 1751266522
transform 1 0 1148 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1751266522
transform -1 0 1212 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1751266522
transform 1 0 1212 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_202
timestamp 1751266522
transform -1 0 1260 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_79
timestamp 1751266522
transform -1 0 1292 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_44
timestamp 1751266522
transform 1 0 1292 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_27
timestamp 1751266522
transform -1 0 1364 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_9
timestamp 1751266522
transform -1 0 1396 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_115
timestamp 1751266522
transform 1 0 1396 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_2_0
timestamp 1751266522
transform 1 0 1428 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1751266522
transform 1 0 1436 0 1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_47
timestamp 1751266522
transform 1 0 1444 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_241
timestamp 1751266522
transform 1 0 1476 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_44
timestamp 1751266522
transform -1 0 1524 0 1 1705
box -2 -3 18 103
use OAI22X1  OAI22X1_6
timestamp 1751266522
transform -1 0 1564 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_2
timestamp 1751266522
transform -1 0 1596 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1751266522
transform 1 0 1596 0 1 1705
box -2 -3 18 103
use BUFX4  BUFX4_240
timestamp 1751266522
transform 1 0 1612 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_17
timestamp 1751266522
transform 1 0 1644 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_19
timestamp 1751266522
transform -1 0 1708 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_20
timestamp 1751266522
transform 1 0 1708 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_33
timestamp 1751266522
transform -1 0 1740 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_34
timestamp 1751266522
transform -1 0 1756 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_136
timestamp 1751266522
transform 1 0 1756 0 1 1705
box -2 -3 26 103
use DFFSR  DFFSR_227
timestamp 1751266522
transform -1 0 1956 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_3_0
timestamp 1751266522
transform 1 0 1956 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1751266522
transform 1 0 1964 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_120
timestamp 1751266522
transform 1 0 1972 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_298
timestamp 1751266522
transform 1 0 1988 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_65
timestamp 1751266522
transform -1 0 2060 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_297
timestamp 1751266522
transform 1 0 2060 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_107
timestamp 1751266522
transform 1 0 2092 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_108
timestamp 1751266522
transform -1 0 2140 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_138
timestamp 1751266522
transform 1 0 2140 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_143
timestamp 1751266522
transform 1 0 2164 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_279
timestamp 1751266522
transform 1 0 2188 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_345
timestamp 1751266522
transform 1 0 2220 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_156
timestamp 1751266522
transform 1 0 2252 0 1 1705
box -2 -3 18 103
use DFFSR  DFFSR_117
timestamp 1751266522
transform -1 0 2444 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_4_0
timestamp 1751266522
transform -1 0 2452 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1751266522
transform -1 0 2460 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_659
timestamp 1751266522
transform -1 0 2492 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1751266522
transform -1 0 2508 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_242
timestamp 1751266522
transform 1 0 2508 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_660
timestamp 1751266522
transform 1 0 2532 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_242
timestamp 1751266522
transform 1 0 2564 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_658
timestamp 1751266522
transform -1 0 2620 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_166
timestamp 1751266522
transform -1 0 2652 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_201
timestamp 1751266522
transform 1 0 2652 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_576
timestamp 1751266522
transform -1 0 2716 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_199
timestamp 1751266522
transform 1 0 2716 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_171
timestamp 1751266522
transform 1 0 2740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_524
timestamp 1751266522
transform 1 0 2772 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_107
timestamp 1751266522
transform -1 0 2844 0 1 1705
box -2 -3 42 103
use INVX1  INVX1_154
timestamp 1751266522
transform -1 0 2860 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_599
timestamp 1751266522
transform -1 0 2892 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_5_0
timestamp 1751266522
transform -1 0 2900 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1751266522
transform -1 0 2908 0 1 1705
box -2 -3 10 103
use DFFSR  DFFSR_172
timestamp 1751266522
transform -1 0 3084 0 1 1705
box -2 -3 178 103
use OAI21X1  OAI21X1_478
timestamp 1751266522
transform 1 0 3084 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_181
timestamp 1751266522
transform -1 0 3140 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_479
timestamp 1751266522
transform 1 0 3140 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_94
timestamp 1751266522
transform 1 0 3172 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_154
timestamp 1751266522
transform -1 0 3244 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_477
timestamp 1751266522
transform -1 0 3276 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_436
timestamp 1751266522
transform 1 0 3276 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_88
timestamp 1751266522
transform 1 0 3308 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_198
timestamp 1751266522
transform 1 0 3348 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_434
timestamp 1751266522
transform -1 0 3404 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_142
timestamp 1751266522
transform -1 0 3436 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_170
timestamp 1751266522
transform 1 0 3436 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_6_0
timestamp 1751266522
transform -1 0 3468 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1751266522
transform -1 0 3476 0 1 1705
box -2 -3 10 103
use BUFX4  BUFX4_252
timestamp 1751266522
transform -1 0 3508 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_153
timestamp 1751266522
transform -1 0 3540 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_155
timestamp 1751266522
transform -1 0 3556 0 1 1705
box -2 -3 18 103
use BUFX4  BUFX4_125
timestamp 1751266522
transform -1 0 3588 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_179
timestamp 1751266522
transform 1 0 3588 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_433
timestamp 1751266522
transform 1 0 3612 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_484
timestamp 1751266522
transform -1 0 3676 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_483
timestamp 1751266522
transform 1 0 3676 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_156
timestamp 1751266522
transform -1 0 3740 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_153
timestamp 1751266522
transform -1 0 3756 0 1 1705
box -2 -3 18 103
use INVX2  INVX2_152
timestamp 1751266522
transform -1 0 3772 0 1 1705
box -2 -3 18 103
use INVX2  INVX2_142
timestamp 1751266522
transform -1 0 3788 0 1 1705
box -2 -3 18 103
use DFFSR  DFFSR_220
timestamp 1751266522
transform -1 0 3964 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_7_0
timestamp 1751266522
transform 1 0 3964 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_7_1
timestamp 1751266522
transform 1 0 3972 0 1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_151
timestamp 1751266522
transform 1 0 3980 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_155
timestamp 1751266522
transform -1 0 4044 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_230
timestamp 1751266522
transform 1 0 4044 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_157
timestamp 1751266522
transform -1 0 4108 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_237
timestamp 1751266522
transform 1 0 4108 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_238
timestamp 1751266522
transform -1 0 4172 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_233
timestamp 1751266522
transform 1 0 4172 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1751266522
transform 1 0 4204 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_207
timestamp 1751266522
transform -1 0 4268 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_158
timestamp 1751266522
transform -1 0 4300 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_211
timestamp 1751266522
transform 1 0 4300 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_58
timestamp 1751266522
transform -1 0 4364 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_142
timestamp 1751266522
transform -1 0 4396 0 1 1705
box -2 -3 34 103
use BUFX2  BUFX2_9
timestamp 1751266522
transform -1 0 28 0 -1 1905
box -2 -3 26 103
use BUFX2  BUFX2_49
timestamp 1751266522
transform -1 0 52 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_132
timestamp 1751266522
transform 1 0 52 0 -1 1905
box -2 -3 34 103
use DFFSR  DFFSR_78
timestamp 1751266522
transform -1 0 260 0 -1 1905
box -2 -3 178 103
use INVX2  INVX2_13
timestamp 1751266522
transform 1 0 260 0 -1 1905
box -2 -3 18 103
use DFFSR  DFFSR_26
timestamp 1751266522
transform -1 0 452 0 -1 1905
box -2 -3 178 103
use FILL  FILL_18_0_0
timestamp 1751266522
transform 1 0 452 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1751266522
transform 1 0 460 0 -1 1905
box -2 -3 10 103
use DFFSR  DFFSR_48
timestamp 1751266522
transform 1 0 468 0 -1 1905
box -2 -3 178 103
use OAI21X1  OAI21X1_56
timestamp 1751266522
transform 1 0 644 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1751266522
transform -1 0 708 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1751266522
transform -1 0 740 0 -1 1905
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1751266522
transform -1 0 772 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1751266522
transform 1 0 772 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_40
timestamp 1751266522
transform -1 0 844 0 -1 1905
box -2 -3 42 103
use OAI22X1  OAI22X1_5
timestamp 1751266522
transform 1 0 844 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_109
timestamp 1751266522
transform 1 0 884 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_1_0
timestamp 1751266522
transform 1 0 916 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1751266522
transform 1 0 924 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_111
timestamp 1751266522
transform 1 0 932 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1751266522
transform -1 0 1004 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_74
timestamp 1751266522
transform 1 0 1004 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_123
timestamp 1751266522
transform 1 0 1036 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_220
timestamp 1751266522
transform 1 0 1068 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_40
timestamp 1751266522
transform -1 0 1132 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1751266522
transform -1 0 1164 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1751266522
transform 1 0 1164 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1751266522
transform 1 0 1196 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1751266522
transform -1 0 1244 0 -1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_4
timestamp 1751266522
transform 1 0 1244 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_3
timestamp 1751266522
transform 1 0 1276 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_80
timestamp 1751266522
transform -1 0 1340 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_600
timestamp 1751266522
transform 1 0 1340 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_64
timestamp 1751266522
transform 1 0 1372 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_85
timestamp 1751266522
transform 1 0 1396 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_2_0
timestamp 1751266522
transform -1 0 1436 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1751266522
transform -1 0 1444 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_77
timestamp 1751266522
transform -1 0 1476 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1751266522
transform -1 0 1508 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_3
timestamp 1751266522
transform 1 0 1508 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_36
timestamp 1751266522
transform -1 0 1556 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_27
timestamp 1751266522
transform -1 0 1572 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_7
timestamp 1751266522
transform 1 0 1572 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1751266522
transform -1 0 1620 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1751266522
transform 1 0 1620 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_18
timestamp 1751266522
transform 1 0 1652 0 -1 1905
box -2 -3 42 103
use OAI22X1  OAI22X1_3
timestamp 1751266522
transform -1 0 1732 0 -1 1905
box -2 -3 42 103
use INVX2  INVX2_24
timestamp 1751266522
transform -1 0 1748 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_2
timestamp 1751266522
transform -1 0 1772 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_35
timestamp 1751266522
transform -1 0 1788 0 -1 1905
box -2 -3 18 103
use DFFSR  DFFSR_121
timestamp 1751266522
transform 1 0 1788 0 -1 1905
box -2 -3 178 103
use FILL  FILL_18_3_0
timestamp 1751266522
transform 1 0 1964 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1751266522
transform 1 0 1972 0 -1 1905
box -2 -3 10 103
use BUFX4  BUFX4_77
timestamp 1751266522
transform 1 0 1980 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_102
timestamp 1751266522
transform 1 0 2012 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_302
timestamp 1751266522
transform 1 0 2028 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_173
timestamp 1751266522
transform -1 0 2092 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_20
timestamp 1751266522
transform -1 0 2140 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_28
timestamp 1751266522
transform -1 0 2188 0 -1 1905
box -2 -3 50 103
use NAND3X1  NAND3X1_274
timestamp 1751266522
transform -1 0 2220 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_220
timestamp 1751266522
transform 1 0 2220 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_29
timestamp 1751266522
transform 1 0 2244 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_646
timestamp 1751266522
transform 1 0 2276 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_645
timestamp 1751266522
transform -1 0 2340 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_236
timestamp 1751266522
transform -1 0 2364 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_239
timestamp 1751266522
transform 1 0 2364 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_121
timestamp 1751266522
transform 1 0 2388 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_644
timestamp 1751266522
transform -1 0 2436 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_4_0
timestamp 1751266522
transform 1 0 2436 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1751266522
transform 1 0 2444 0 -1 1905
box -2 -3 10 103
use INVX2  INVX2_143
timestamp 1751266522
transform 1 0 2452 0 -1 1905
box -2 -3 18 103
use BUFX4  BUFX4_18
timestamp 1751266522
transform 1 0 2468 0 -1 1905
box -2 -3 34 103
use DFFSR  DFFSR_185
timestamp 1751266522
transform -1 0 2676 0 -1 1905
box -2 -3 178 103
use AOI21X1  AOI21X1_190
timestamp 1751266522
transform -1 0 2708 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_563
timestamp 1751266522
transform -1 0 2740 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_211
timestamp 1751266522
transform 1 0 2740 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_147
timestamp 1751266522
transform -1 0 2796 0 -1 1905
box -2 -3 34 103
use INVX2  INVX2_102
timestamp 1751266522
transform 1 0 2796 0 -1 1905
box -2 -3 18 103
use CLKBUF1  CLKBUF1_21
timestamp 1751266522
transform 1 0 2812 0 -1 1905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_65
timestamp 1751266522
transform -1 0 2956 0 -1 1905
box -2 -3 74 103
use FILL  FILL_18_5_0
timestamp 1751266522
transform 1 0 2956 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1751266522
transform 1 0 2964 0 -1 1905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_9
timestamp 1751266522
transform 1 0 2972 0 -1 1905
box -2 -3 74 103
use BUFX4  BUFX4_41
timestamp 1751266522
transform 1 0 3044 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_98
timestamp 1751266522
transform 1 0 3076 0 -1 1905
box -2 -3 42 103
use AOI21X1  AOI21X1_158
timestamp 1751266522
transform 1 0 3116 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_489
timestamp 1751266522
transform 1 0 3148 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1751266522
transform -1 0 3212 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_490
timestamp 1751266522
transform 1 0 3212 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_232
timestamp 1751266522
transform -1 0 3276 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_398
timestamp 1751266522
transform -1 0 3308 0 -1 1905
box -2 -3 34 103
use INVX2  INVX2_100
timestamp 1751266522
transform 1 0 3308 0 -1 1905
box -2 -3 18 103
use DFFSR  DFFSR_217
timestamp 1751266522
transform -1 0 3500 0 -1 1905
box -2 -3 178 103
use FILL  FILL_18_6_0
timestamp 1751266522
transform 1 0 3500 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1751266522
transform 1 0 3508 0 -1 1905
box -2 -3 10 103
use AOI22X1  AOI22X1_55
timestamp 1751266522
transform 1 0 3516 0 -1 1905
box -2 -3 42 103
use BUFX4  BUFX4_247
timestamp 1751266522
transform -1 0 3588 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_397
timestamp 1751266522
transform 1 0 3588 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_124
timestamp 1751266522
transform -1 0 3652 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_394
timestamp 1751266522
transform -1 0 3684 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_121
timestamp 1751266522
transform 1 0 3684 0 -1 1905
box -2 -3 34 103
use INVX2  INVX2_158
timestamp 1751266522
transform 1 0 3716 0 -1 1905
box -2 -3 18 103
use AOI22X1  AOI22X1_53
timestamp 1751266522
transform 1 0 3732 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_393
timestamp 1751266522
transform 1 0 3772 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_120
timestamp 1751266522
transform -1 0 3836 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_189
timestamp 1751266522
transform -1 0 3860 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_152
timestamp 1751266522
transform -1 0 3884 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_159
timestamp 1751266522
transform -1 0 3900 0 -1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_154
timestamp 1751266522
transform 1 0 3900 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_150
timestamp 1751266522
transform 1 0 3932 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_7_0
timestamp 1751266522
transform -1 0 3972 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_7_1
timestamp 1751266522
transform -1 0 3980 0 -1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_152
timestamp 1751266522
transform -1 0 4012 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_156
timestamp 1751266522
transform 1 0 4012 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_74
timestamp 1751266522
transform 1 0 4044 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_144
timestamp 1751266522
transform -1 0 4092 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_132
timestamp 1751266522
transform -1 0 4108 0 -1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_236
timestamp 1751266522
transform 1 0 4108 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_234
timestamp 1751266522
transform 1 0 4140 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_235
timestamp 1751266522
transform -1 0 4204 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_75
timestamp 1751266522
transform -1 0 4236 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_6
timestamp 1751266522
transform 1 0 4236 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_49
timestamp 1751266522
transform -1 0 4300 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_86
timestamp 1751266522
transform -1 0 4316 0 -1 1905
box -2 -3 18 103
use INVX2  INVX2_66
timestamp 1751266522
transform -1 0 4332 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_215
timestamp 1751266522
transform -1 0 4364 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_64
timestamp 1751266522
transform -1 0 4388 0 -1 1905
box -2 -3 26 103
use FILL  FILL_19_1
timestamp 1751266522
transform -1 0 4396 0 -1 1905
box -2 -3 10 103
use BUFX2  BUFX2_8
timestamp 1751266522
transform -1 0 28 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_28
timestamp 1751266522
transform -1 0 52 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_131
timestamp 1751266522
transform 1 0 52 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_151
timestamp 1751266522
transform 1 0 84 0 1 1905
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1751266522
transform -1 0 140 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_13
timestamp 1751266522
transform -1 0 164 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_129
timestamp 1751266522
transform 1 0 164 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_136
timestamp 1751266522
transform 1 0 196 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_15
timestamp 1751266522
transform 1 0 228 0 1 1905
box -2 -3 18 103
use DFFSR  DFFSR_6
timestamp 1751266522
transform -1 0 420 0 1 1905
box -2 -3 178 103
use FILL  FILL_19_0_0
timestamp 1751266522
transform -1 0 428 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1751266522
transform -1 0 436 0 1 1905
box -2 -3 10 103
use DFFSR  DFFSR_11
timestamp 1751266522
transform -1 0 612 0 1 1905
box -2 -3 178 103
use INVX2  INVX2_4
timestamp 1751266522
transform 1 0 612 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_60
timestamp 1751266522
transform 1 0 628 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_38
timestamp 1751266522
transform 1 0 660 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_32
timestamp 1751266522
transform -1 0 724 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1751266522
transform 1 0 724 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_57
timestamp 1751266522
transform 1 0 756 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1751266522
transform -1 0 820 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1751266522
transform 1 0 820 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_128
timestamp 1751266522
transform -1 0 884 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_40
timestamp 1751266522
transform 1 0 884 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_1_0
timestamp 1751266522
transform 1 0 900 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1751266522
transform 1 0 908 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_112
timestamp 1751266522
transform 1 0 916 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1751266522
transform 1 0 948 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_59
timestamp 1751266522
transform -1 0 1012 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_66
timestamp 1751266522
transform 1 0 1012 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_67
timestamp 1751266522
transform -1 0 1076 0 1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_16
timestamp 1751266522
transform -1 0 1116 0 1 1905
box -2 -3 42 103
use NOR2X1  NOR2X1_15
timestamp 1751266522
transform 1 0 1116 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_48
timestamp 1751266522
transform -1 0 1164 0 1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_49
timestamp 1751266522
transform 1 0 1164 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_8
timestamp 1751266522
transform 1 0 1196 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1751266522
transform 1 0 1228 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_25
timestamp 1751266522
transform -1 0 1276 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_4
timestamp 1751266522
transform 1 0 1276 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1751266522
transform 1 0 1292 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1751266522
transform 1 0 1324 0 1 1905
box -2 -3 26 103
use OAI22X1  OAI22X1_42
timestamp 1751266522
transform -1 0 1388 0 1 1905
box -2 -3 42 103
use AOI21X1  AOI21X1_14
timestamp 1751266522
transform -1 0 1420 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1751266522
transform 1 0 1420 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1751266522
transform 1 0 1428 0 1 1905
box -2 -3 10 103
use AOI22X1  AOI22X1_28
timestamp 1751266522
transform 1 0 1436 0 1 1905
box -2 -3 42 103
use NAND3X1  NAND3X1_43
timestamp 1751266522
transform 1 0 1476 0 1 1905
box -2 -3 34 103
use DFFSR  DFFSR_34
timestamp 1751266522
transform 1 0 1508 0 1 1905
box -2 -3 178 103
use AOI21X1  AOI21X1_1
timestamp 1751266522
transform 1 0 1684 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1751266522
transform -1 0 1740 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_35
timestamp 1751266522
transform 1 0 1740 0 1 1905
box -2 -3 26 103
use OAI22X1  OAI22X1_41
timestamp 1751266522
transform 1 0 1764 0 1 1905
box -2 -3 42 103
use INVX8  INVX8_20
timestamp 1751266522
transform 1 0 1804 0 1 1905
box -2 -3 42 103
use BUFX4  BUFX4_91
timestamp 1751266522
transform 1 0 1844 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_90
timestamp 1751266522
transform 1 0 1876 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_140
timestamp 1751266522
transform 1 0 1908 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_3_0
timestamp 1751266522
transform -1 0 1940 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1751266522
transform -1 0 1948 0 1 1905
box -2 -3 10 103
use INVX1  INVX1_57
timestamp 1751266522
transform -1 0 1964 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_59
timestamp 1751266522
transform -1 0 1980 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_185
timestamp 1751266522
transform -1 0 2004 0 1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_27
timestamp 1751266522
transform -1 0 2044 0 1 1905
box -2 -3 42 103
use BUFX4  BUFX4_168
timestamp 1751266522
transform -1 0 2076 0 1 1905
box -2 -3 34 103
use DFFSR  DFFSR_124
timestamp 1751266522
transform -1 0 2252 0 1 1905
box -2 -3 178 103
use NOR2X1  NOR2X1_215
timestamp 1751266522
transform 1 0 2252 0 1 1905
box -2 -3 26 103
use DFFSR  DFFSR_156
timestamp 1751266522
transform -1 0 2452 0 1 1905
box -2 -3 178 103
use FILL  FILL_19_4_0
timestamp 1751266522
transform 1 0 2452 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1751266522
transform 1 0 2460 0 1 1905
box -2 -3 10 103
use OAI22X1  OAI22X1_116
timestamp 1751266522
transform 1 0 2468 0 1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_565
timestamp 1751266522
transform -1 0 2540 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_564
timestamp 1751266522
transform -1 0 2572 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_101
timestamp 1751266522
transform 1 0 2572 0 1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_12
timestamp 1751266522
transform 1 0 2588 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_180
timestamp 1751266522
transform -1 0 2660 0 1 1905
box -2 -3 26 103
use DFFSR  DFFSR_193
timestamp 1751266522
transform -1 0 2836 0 1 1905
box -2 -3 178 103
use DFFSR  DFFSR_241
timestamp 1751266522
transform -1 0 3012 0 1 1905
box -2 -3 178 103
use FILL  FILL_19_5_0
timestamp 1751266522
transform 1 0 3012 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1751266522
transform 1 0 3020 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_469
timestamp 1751266522
transform 1 0 3028 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_353
timestamp 1751266522
transform 1 0 3060 0 1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_91
timestamp 1751266522
transform 1 0 3092 0 1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_470
timestamp 1751266522
transform -1 0 3164 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_151
timestamp 1751266522
transform -1 0 3196 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_468
timestamp 1751266522
transform -1 0 3228 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_174
timestamp 1751266522
transform -1 0 3252 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1751266522
transform 1 0 3252 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_231
timestamp 1751266522
transform -1 0 3316 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_82
timestamp 1751266522
transform -1 0 3348 0 1 1905
box -2 -3 34 103
use INVX8  INVX8_18
timestamp 1751266522
transform 1 0 3348 0 1 1905
box -2 -3 42 103
use AOI22X1  AOI22X1_37
timestamp 1751266522
transform 1 0 3388 0 1 1905
box -2 -3 42 103
use AOI21X1  AOI21X1_125
timestamp 1751266522
transform 1 0 3428 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_6_0
timestamp 1751266522
transform -1 0 3468 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1751266522
transform -1 0 3476 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_243
timestamp 1751266522
transform -1 0 3508 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_413
timestamp 1751266522
transform -1 0 3540 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_352
timestamp 1751266522
transform 1 0 3540 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_82
timestamp 1751266522
transform -1 0 3604 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1751266522
transform -1 0 3628 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_149
timestamp 1751266522
transform -1 0 3652 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_151
timestamp 1751266522
transform -1 0 3676 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_147
timestamp 1751266522
transform 1 0 3676 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_148
timestamp 1751266522
transform 1 0 3700 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_267
timestamp 1751266522
transform 1 0 3724 0 1 1905
box -2 -3 34 103
use DFFSR  DFFSR_225
timestamp 1751266522
transform -1 0 3932 0 1 1905
box -2 -3 178 103
use NOR2X1  NOR2X1_85
timestamp 1751266522
transform 1 0 3932 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_137
timestamp 1751266522
transform -1 0 3980 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_7_0
timestamp 1751266522
transform 1 0 3980 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_7_1
timestamp 1751266522
transform 1 0 3988 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_134
timestamp 1751266522
transform 1 0 3996 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_135
timestamp 1751266522
transform 1 0 4020 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_133
timestamp 1751266522
transform 1 0 4036 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_94
timestamp 1751266522
transform 1 0 4052 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_111
timestamp 1751266522
transform 1 0 4076 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_63
timestamp 1751266522
transform 1 0 4100 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_104
timestamp 1751266522
transform -1 0 4164 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1751266522
transform 1 0 4164 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_231
timestamp 1751266522
transform -1 0 4228 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_251
timestamp 1751266522
transform -1 0 4260 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_127
timestamp 1751266522
transform -1 0 4292 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_63
timestamp 1751266522
transform 1 0 4292 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_92
timestamp 1751266522
transform 1 0 4316 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_32
timestamp 1751266522
transform -1 0 4372 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1751266522
transform 1 0 4372 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1751266522
transform 1 0 4380 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_3
timestamp 1751266522
transform 1 0 4388 0 1 1905
box -2 -3 10 103
use BUFX2  BUFX2_4
timestamp 1751266522
transform -1 0 28 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_127
timestamp 1751266522
transform -1 0 60 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1751266522
transform 1 0 60 0 -1 2105
box -2 -3 18 103
use DFFSR  DFFSR_2
timestamp 1751266522
transform -1 0 252 0 -1 2105
box -2 -3 178 103
use DFFSR  DFFSR_62
timestamp 1751266522
transform 1 0 252 0 -1 2105
box -2 -3 178 103
use FILL  FILL_20_0_0
timestamp 1751266522
transform 1 0 428 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1751266522
transform 1 0 436 0 -1 2105
box -2 -3 10 103
use INVX2  INVX2_38
timestamp 1751266522
transform 1 0 444 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_108
timestamp 1751266522
transform 1 0 460 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1751266522
transform 1 0 492 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_36
timestamp 1751266522
transform -1 0 540 0 -1 2105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_43
timestamp 1751266522
transform -1 0 612 0 -1 2105
box -2 -3 74 103
use INVX2  INVX2_39
timestamp 1751266522
transform 1 0 612 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_1
timestamp 1751266522
transform -1 0 652 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_110
timestamp 1751266522
transform 1 0 652 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1751266522
transform -1 0 716 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_30
timestamp 1751266522
transform 1 0 716 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_59
timestamp 1751266522
transform 1 0 732 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1751266522
transform -1 0 796 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1751266522
transform 1 0 796 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_130
timestamp 1751266522
transform -1 0 860 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1751266522
transform 1 0 860 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_1_0
timestamp 1751266522
transform -1 0 900 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1751266522
transform -1 0 908 0 -1 2105
box -2 -3 10 103
use BUFX4  BUFX4_131
timestamp 1751266522
transform -1 0 940 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_37
timestamp 1751266522
transform 1 0 940 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_92
timestamp 1751266522
transform -1 0 1004 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_32
timestamp 1751266522
transform 1 0 1004 0 -1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_124
timestamp 1751266522
transform 1 0 1044 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_210
timestamp 1751266522
transform 1 0 1076 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1751266522
transform -1 0 1140 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_48
timestamp 1751266522
transform 1 0 1140 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1751266522
transform -1 0 1204 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_38
timestamp 1751266522
transform 1 0 1204 0 -1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_83
timestamp 1751266522
transform -1 0 1412 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_2_0
timestamp 1751266522
transform 1 0 1412 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1751266522
transform 1 0 1420 0 -1 2105
box -2 -3 10 103
use BUFX4  BUFX4_117
timestamp 1751266522
transform 1 0 1428 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_78
timestamp 1751266522
transform 1 0 1460 0 -1 2105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_25
timestamp 1751266522
transform 1 0 1492 0 -1 2105
box -2 -3 74 103
use BUFX2  BUFX2_75
timestamp 1751266522
transform 1 0 1564 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_28
timestamp 1751266522
transform 1 0 1588 0 -1 2105
box -2 -3 18 103
use INVX2  INVX2_23
timestamp 1751266522
transform 1 0 1604 0 -1 2105
box -2 -3 18 103
use DFFSR  DFFSR_116
timestamp 1751266522
transform -1 0 1796 0 -1 2105
box -2 -3 178 103
use INVX1  INVX1_58
timestamp 1751266522
transform -1 0 1812 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_268
timestamp 1751266522
transform -1 0 1844 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_267
timestamp 1751266522
transform 1 0 1844 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_54
timestamp 1751266522
transform -1 0 1916 0 -1 2105
box -2 -3 42 103
use FILL  FILL_20_3_0
timestamp 1751266522
transform -1 0 1924 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1751266522
transform -1 0 1932 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_291
timestamp 1751266522
transform -1 0 1964 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_83
timestamp 1751266522
transform 1 0 1964 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_84
timestamp 1751266522
transform -1 0 2012 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_265
timestamp 1751266522
transform 1 0 2012 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_82
timestamp 1751266522
transform 1 0 2044 0 -1 2105
box -2 -3 26 103
use OAI22X1  OAI22X1_53
timestamp 1751266522
transform -1 0 2108 0 -1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_81
timestamp 1751266522
transform -1 0 2132 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_264
timestamp 1751266522
transform -1 0 2164 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_276
timestamp 1751266522
transform 1 0 2164 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_177
timestamp 1751266522
transform -1 0 2372 0 -1 2105
box -2 -3 178 103
use NOR2X1  NOR2X1_231
timestamp 1751266522
transform -1 0 2396 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_90
timestamp 1751266522
transform 1 0 2396 0 -1 2105
box -2 -3 18 103
use OAI22X1  OAI22X1_103
timestamp 1751266522
transform 1 0 2412 0 -1 2105
box -2 -3 42 103
use FILL  FILL_20_4_0
timestamp 1751266522
transform 1 0 2452 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1751266522
transform 1 0 2460 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_631
timestamp 1751266522
transform 1 0 2468 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_632
timestamp 1751266522
transform 1 0 2500 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_129
timestamp 1751266522
transform -1 0 2708 0 -1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_512
timestamp 1751266522
transform -1 0 2740 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_511
timestamp 1751266522
transform 1 0 2740 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_235
timestamp 1751266522
transform 1 0 2772 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_630
timestamp 1751266522
transform 1 0 2796 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_112
timestamp 1751266522
transform -1 0 2868 0 -1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_551
timestamp 1751266522
transform -1 0 2900 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_550
timestamp 1751266522
transform 1 0 2900 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_86
timestamp 1751266522
transform 1 0 2932 0 -1 2105
box -2 -3 18 103
use FILL  FILL_20_5_0
timestamp 1751266522
transform 1 0 2948 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1751266522
transform 1 0 2956 0 -1 2105
box -2 -3 10 103
use INVX2  INVX2_87
timestamp 1751266522
transform 1 0 2964 0 -1 2105
box -2 -3 18 103
use INVX2  INVX2_88
timestamp 1751266522
transform -1 0 2996 0 -1 2105
box -2 -3 18 103
use DFFSR  DFFSR_209
timestamp 1751266522
transform -1 0 3172 0 -1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_415
timestamp 1751266522
transform -1 0 3204 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_416
timestamp 1751266522
transform 1 0 3204 0 -1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_83
timestamp 1751266522
transform 1 0 3236 0 -1 2105
box -2 -3 42 103
use AOI21X1  AOI21X1_137
timestamp 1751266522
transform 1 0 3276 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_414
timestamp 1751266522
transform -1 0 3340 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1751266522
transform -1 0 3364 0 -1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_10
timestamp 1751266522
transform 1 0 3364 0 -1 2105
box -2 -3 50 103
use OAI21X1  OAI21X1_357
timestamp 1751266522
transform -1 0 3444 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_87
timestamp 1751266522
transform 1 0 3444 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_6_0
timestamp 1751266522
transform -1 0 3484 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1751266522
transform -1 0 3492 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_383
timestamp 1751266522
transform -1 0 3524 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_111
timestamp 1751266522
transform -1 0 3556 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1751266522
transform -1 0 3580 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_183
timestamp 1751266522
transform -1 0 3604 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_421
timestamp 1751266522
transform -1 0 3636 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_85
timestamp 1751266522
transform -1 0 3652 0 -1 2105
box -2 -3 18 103
use BUFX4  BUFX4_250
timestamp 1751266522
transform 1 0 3652 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_179
timestamp 1751266522
transform 1 0 3684 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_110
timestamp 1751266522
transform 1 0 3708 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_382
timestamp 1751266522
transform -1 0 3772 0 -1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_49
timestamp 1751266522
transform -1 0 3812 0 -1 2105
box -2 -3 42 103
use BUFX4  BUFX4_156
timestamp 1751266522
transform 1 0 3812 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_9
timestamp 1751266522
transform 1 0 3844 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_105
timestamp 1751266522
transform 1 0 3892 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_72
timestamp 1751266522
transform -1 0 3940 0 -1 2105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_54
timestamp 1751266522
transform -1 0 4012 0 -1 2105
box -2 -3 74 103
use FILL  FILL_20_7_0
timestamp 1751266522
transform 1 0 4012 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_7_1
timestamp 1751266522
transform 1 0 4020 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_107
timestamp 1751266522
transform 1 0 4028 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_43
timestamp 1751266522
transform 1 0 4052 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_214
timestamp 1751266522
transform -1 0 4116 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_214
timestamp 1751266522
transform 1 0 4116 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_207
timestamp 1751266522
transform -1 0 4180 0 -1 2105
box -2 -3 34 103
use NOR3X1  NOR3X1_4
timestamp 1751266522
transform 1 0 4180 0 -1 2105
box -2 -3 66 103
use INVX1  INVX1_107
timestamp 1751266522
transform 1 0 4244 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_160
timestamp 1751266522
transform 1 0 4260 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_159
timestamp 1751266522
transform 1 0 4292 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_223
timestamp 1751266522
transform 1 0 4324 0 -1 2105
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1751266522
transform 1 0 4356 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_90
timestamp 1751266522
transform -1 0 4396 0 -1 2105
box -2 -3 18 103
use BUFX2  BUFX2_31
timestamp 1751266522
transform -1 0 28 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_61
timestamp 1751266522
transform -1 0 52 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_15
timestamp 1751266522
transform -1 0 76 0 1 2105
box -2 -3 26 103
use DFFSR  DFFSR_90
timestamp 1751266522
transform -1 0 252 0 1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_138
timestamp 1751266522
transform -1 0 284 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1751266522
transform 1 0 284 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1751266522
transform 1 0 316 0 1 2105
box -2 -3 18 103
use FILL  FILL_21_0_0
timestamp 1751266522
transform 1 0 332 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1751266522
transform 1 0 340 0 1 2105
box -2 -3 10 103
use DFFSR  DFFSR_60
timestamp 1751266522
transform 1 0 348 0 1 2105
box -2 -3 178 103
use DFFSR  DFFSR_47
timestamp 1751266522
transform -1 0 700 0 1 2105
box -2 -3 178 103
use BUFX4  BUFX4_200
timestamp 1751266522
transform 1 0 700 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_63
timestamp 1751266522
transform -1 0 764 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_42
timestamp 1751266522
transform 1 0 764 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_65
timestamp 1751266522
transform 1 0 796 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1751266522
transform 1 0 828 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1751266522
transform 1 0 860 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_1_0
timestamp 1751266522
transform 1 0 892 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1751266522
transform 1 0 900 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_41
timestamp 1751266522
transform 1 0 908 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1751266522
transform 1 0 940 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_202
timestamp 1751266522
transform -1 0 1004 0 1 2105
box -2 -3 34 103
use OAI22X1  OAI22X1_38
timestamp 1751266522
transform 1 0 1004 0 1 2105
box -2 -3 42 103
use OAI22X1  OAI22X1_35
timestamp 1751266522
transform -1 0 1084 0 1 2105
box -2 -3 42 103
use BUFX4  BUFX4_196
timestamp 1751266522
transform -1 0 1116 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1751266522
transform -1 0 1140 0 1 2105
box -2 -3 26 103
use DFFSR  DFFSR_29
timestamp 1751266522
transform -1 0 1316 0 1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_10
timestamp 1751266522
transform 1 0 1316 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1751266522
transform 1 0 1348 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1751266522
transform -1 0 1396 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_9
timestamp 1751266522
transform 1 0 1396 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_2_0
timestamp 1751266522
transform 1 0 1428 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1751266522
transform 1 0 1436 0 1 2105
box -2 -3 10 103
use DFFSR  DFFSR_37
timestamp 1751266522
transform 1 0 1444 0 1 2105
box -2 -3 178 103
use AOI22X1  AOI22X1_26
timestamp 1751266522
transform 1 0 1620 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_20
timestamp 1751266522
transform 1 0 1660 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_24
timestamp 1751266522
transform 1 0 1700 0 1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_18
timestamp 1751266522
transform 1 0 1740 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_83
timestamp 1751266522
transform 1 0 1764 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_81
timestamp 1751266522
transform 1 0 1796 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_86
timestamp 1751266522
transform -1 0 1860 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_89
timestamp 1751266522
transform 1 0 1860 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_266
timestamp 1751266522
transform 1 0 1892 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_3_0
timestamp 1751266522
transform -1 0 1932 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1751266522
transform -1 0 1940 0 1 2105
box -2 -3 10 103
use OAI22X1  OAI22X1_61
timestamp 1751266522
transform -1 0 1980 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_288
timestamp 1751266522
transform -1 0 2012 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_287
timestamp 1751266522
transform -1 0 2044 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_318
timestamp 1751266522
transform -1 0 2076 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1751266522
transform 1 0 2076 0 1 2105
box -2 -3 26 103
use OAI22X1  OAI22X1_73
timestamp 1751266522
transform -1 0 2140 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_319
timestamp 1751266522
transform -1 0 2172 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_322
timestamp 1751266522
transform 1 0 2172 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_53
timestamp 1751266522
transform -1 0 2220 0 1 2105
box -2 -3 18 103
use BUFX4  BUFX4_225
timestamp 1751266522
transform -1 0 2252 0 1 2105
box -2 -3 34 103
use INVX8  INVX8_22
timestamp 1751266522
transform 1 0 2252 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_347
timestamp 1751266522
transform 1 0 2292 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_584
timestamp 1751266522
transform 1 0 2324 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_162
timestamp 1751266522
transform 1 0 2356 0 1 2105
box -2 -3 34 103
use AND2X2  AND2X2_25
timestamp 1751266522
transform 1 0 2388 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_510
timestamp 1751266522
transform -1 0 2452 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_4_0
timestamp 1751266522
transform -1 0 2460 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1751266522
transform -1 0 2468 0 1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_165
timestamp 1751266522
transform -1 0 2500 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_190
timestamp 1751266522
transform 1 0 2500 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_150
timestamp 1751266522
transform -1 0 2540 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_207
timestamp 1751266522
transform -1 0 2564 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_155
timestamp 1751266522
transform -1 0 2588 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_11
timestamp 1751266522
transform 1 0 2588 0 1 2105
box -2 -3 50 103
use INVX2  INVX2_89
timestamp 1751266522
transform 1 0 2636 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_549
timestamp 1751266522
transform 1 0 2652 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_184
timestamp 1751266522
transform 1 0 2684 0 1 2105
box -2 -3 34 103
use DFFSR  DFFSR_223
timestamp 1751266522
transform -1 0 2892 0 1 2105
box -2 -3 178 103
use INVX2  INVX2_56
timestamp 1751266522
transform 1 0 2892 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_387
timestamp 1751266522
transform -1 0 2940 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_5_0
timestamp 1751266522
transform 1 0 2940 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1751266522
transform 1 0 2948 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_154
timestamp 1751266522
transform 1 0 2956 0 1 2105
box -2 -3 34 103
use DFFSR  DFFSR_239
timestamp 1751266522
transform -1 0 3164 0 1 2105
box -2 -3 178 103
use NOR2X1  NOR2X1_189
timestamp 1751266522
transform 1 0 3164 0 1 2105
box -2 -3 26 103
use INVX2  INVX2_57
timestamp 1751266522
transform 1 0 3188 0 1 2105
box -2 -3 18 103
use AOI21X1  AOI21X1_115
timestamp 1751266522
transform 1 0 3204 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_51
timestamp 1751266522
transform 1 0 3236 0 1 2105
box -2 -3 42 103
use AOI21X1  AOI21X1_119
timestamp 1751266522
transform 1 0 3276 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_39
timestamp 1751266522
transform 1 0 3308 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_356
timestamp 1751266522
transform 1 0 3348 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_86
timestamp 1751266522
transform 1 0 3380 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_386
timestamp 1751266522
transform 1 0 3412 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1751266522
transform -1 0 3476 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_6_0
timestamp 1751266522
transform 1 0 3476 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1751266522
transform 1 0 3484 0 1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_4
timestamp 1751266522
transform 1 0 3492 0 1 2105
box -2 -3 50 103
use BUFX4  BUFX4_263
timestamp 1751266522
transform -1 0 3572 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1751266522
transform 1 0 3572 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_264
timestamp 1751266522
transform -1 0 3636 0 1 2105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_60
timestamp 1751266522
transform 1 0 3636 0 1 2105
box -2 -3 74 103
use NAND2X1  NAND2X1_106
timestamp 1751266522
transform 1 0 3708 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_97
timestamp 1751266522
transform 1 0 3732 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_100
timestamp 1751266522
transform 1 0 3756 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_99
timestamp 1751266522
transform 1 0 3780 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1751266522
transform 1 0 3804 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1751266522
transform 1 0 3836 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1751266522
transform 1 0 3868 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_84
timestamp 1751266522
transform 1 0 3892 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1751266522
transform 1 0 3924 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_55
timestamp 1751266522
transform -1 0 3972 0 1 2105
box -2 -3 18 103
use FILL  FILL_21_7_0
timestamp 1751266522
transform -1 0 3980 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_7_1
timestamp 1751266522
transform -1 0 3988 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_66
timestamp 1751266522
transform -1 0 4020 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_203
timestamp 1751266522
transform -1 0 4052 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_41
timestamp 1751266522
transform 1 0 4052 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_456
timestamp 1751266522
transform -1 0 4116 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1751266522
transform 1 0 4116 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_192
timestamp 1751266522
transform 1 0 4140 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_53
timestamp 1751266522
transform 1 0 4172 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_83
timestamp 1751266522
transform 1 0 4196 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_193
timestamp 1751266522
transform -1 0 4244 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_213
timestamp 1751266522
transform 1 0 4244 0 1 2105
box -2 -3 34 103
use XOR2X1  XOR2X1_5
timestamp 1751266522
transform 1 0 4276 0 1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_7
timestamp 1751266522
transform -1 0 4388 0 1 2105
box -2 -3 58 103
use FILL  FILL_22_1
timestamp 1751266522
transform 1 0 4388 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_67
timestamp 1751266522
transform -1 0 28 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_2
timestamp 1751266522
transform 1 0 28 0 -1 2305
box -2 -3 34 103
use BUFX2  BUFX2_48
timestamp 1751266522
transform -1 0 84 0 -1 2305
box -2 -3 26 103
use DFFSR  DFFSR_77
timestamp 1751266522
transform -1 0 260 0 -1 2305
box -2 -3 178 103
use DFFSR  DFFSR_13
timestamp 1751266522
transform -1 0 436 0 -1 2305
box -2 -3 178 103
use FILL  FILL_22_0_0
timestamp 1751266522
transform 1 0 436 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1751266522
transform 1 0 444 0 -1 2305
box -2 -3 10 103
use DFFSR  DFFSR_40
timestamp 1751266522
transform 1 0 452 0 -1 2305
box -2 -3 178 103
use INVX2  INVX2_34
timestamp 1751266522
transform 1 0 628 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_100
timestamp 1751266522
transform 1 0 644 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1751266522
transform 1 0 676 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_44
timestamp 1751266522
transform 1 0 708 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_116
timestamp 1751266522
transform 1 0 724 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1751266522
transform 1 0 756 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1751266522
transform -1 0 820 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1751266522
transform 1 0 820 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1751266522
transform -1 0 884 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1751266522
transform -1 0 916 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_1_0
timestamp 1751266522
transform -1 0 924 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1751266522
transform -1 0 932 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_101
timestamp 1751266522
transform -1 0 964 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_45
timestamp 1751266522
transform -1 0 980 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_122
timestamp 1751266522
transform 1 0 980 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1751266522
transform 1 0 1012 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_47
timestamp 1751266522
transform -1 0 1060 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1751266522
transform -1 0 1092 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_75
timestamp 1751266522
transform -1 0 1124 0 -1 2305
box -2 -3 34 103
use DFFSR  DFFSR_35
timestamp 1751266522
transform 1 0 1124 0 -1 2305
box -2 -3 178 103
use NAND2X1  NAND2X1_19
timestamp 1751266522
transform 1 0 1300 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_46
timestamp 1751266522
transform -1 0 1356 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_2_0
timestamp 1751266522
transform 1 0 1356 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1751266522
transform 1 0 1364 0 -1 2305
box -2 -3 10 103
use DFFSR  DFFSR_33
timestamp 1751266522
transform 1 0 1372 0 -1 2305
box -2 -3 178 103
use NOR2X1  NOR2X1_13
timestamp 1751266522
transform 1 0 1548 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_46
timestamp 1751266522
transform -1 0 1596 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1751266522
transform 1 0 1596 0 -1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_36
timestamp 1751266522
transform -1 0 1668 0 -1 2305
box -2 -3 42 103
use OAI22X1  OAI22X1_34
timestamp 1751266522
transform 1 0 1668 0 -1 2305
box -2 -3 42 103
use INVX1  INVX1_52
timestamp 1751266522
transform -1 0 1724 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_87
timestamp 1751266522
transform -1 0 1756 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1751266522
transform -1 0 1780 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_38
timestamp 1751266522
transform 1 0 1780 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_99
timestamp 1751266522
transform 1 0 1812 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_100
timestamp 1751266522
transform -1 0 1860 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_91
timestamp 1751266522
transform -1 0 1884 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_275
timestamp 1751266522
transform 1 0 1884 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_3_0
timestamp 1751266522
transform -1 0 1924 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1751266522
transform -1 0 1932 0 -1 2305
box -2 -3 10 103
use OAI22X1  OAI22X1_57
timestamp 1751266522
transform -1 0 1972 0 -1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_90
timestamp 1751266522
transform -1 0 1996 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_274
timestamp 1751266522
transform 1 0 1996 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_51
timestamp 1751266522
transform -1 0 2044 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_278
timestamp 1751266522
transform 1 0 2044 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_124
timestamp 1751266522
transform -1 0 2100 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_125
timestamp 1751266522
transform -1 0 2124 0 -1 2305
box -2 -3 26 103
use DFFSR  DFFSR_143
timestamp 1751266522
transform -1 0 2300 0 -1 2305
box -2 -3 178 103
use AND2X2  AND2X2_26
timestamp 1751266522
transform 1 0 2300 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_233
timestamp 1751266522
transform 1 0 2332 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_636
timestamp 1751266522
transform 1 0 2356 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_217
timestamp 1751266522
transform -1 0 2412 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_21
timestamp 1751266522
transform 1 0 2412 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_4_0
timestamp 1751266522
transform 1 0 2444 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1751266522
transform 1 0 2452 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_592
timestamp 1751266522
transform 1 0 2460 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_593
timestamp 1751266522
transform 1 0 2492 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_224
timestamp 1751266522
transform 1 0 2524 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_93
timestamp 1751266522
transform 1 0 2548 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_590
timestamp 1751266522
transform -1 0 2596 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_3
timestamp 1751266522
transform 1 0 2596 0 -1 2305
box -2 -3 50 103
use DFFSR  DFFSR_161
timestamp 1751266522
transform -1 0 2820 0 -1 2305
box -2 -3 178 103
use INVX2  INVX2_84
timestamp 1751266522
transform 1 0 2820 0 -1 2305
box -2 -3 18 103
use DFFSR  DFFSR_237
timestamp 1751266522
transform -1 0 3012 0 -1 2305
box -2 -3 178 103
use FILL  FILL_22_5_0
timestamp 1751266522
transform -1 0 3020 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1751266522
transform -1 0 3028 0 -1 2305
box -2 -3 10 103
use DFFSR  DFFSR_221
timestamp 1751266522
transform -1 0 3204 0 -1 2305
box -2 -3 178 103
use AOI22X1  AOI22X1_41
timestamp 1751266522
transform 1 0 3204 0 -1 2305
box -2 -3 42 103
use INVX2  INVX2_83
timestamp 1751266522
transform 1 0 3244 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_392
timestamp 1751266522
transform -1 0 3292 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_52
timestamp 1751266522
transform 1 0 3292 0 -1 2305
box -2 -3 42 103
use INVX2  INVX2_128
timestamp 1751266522
transform 1 0 3332 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_8
timestamp 1751266522
transform 1 0 3348 0 -1 2305
box -2 -3 50 103
use AOI21X1  AOI21X1_90
timestamp 1751266522
transform 1 0 3396 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_360
timestamp 1751266522
transform -1 0 3460 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_6_0
timestamp 1751266522
transform 1 0 3460 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1751266522
transform 1 0 3468 0 -1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_118
timestamp 1751266522
transform 1 0 3476 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_391
timestamp 1751266522
transform -1 0 3540 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1751266522
transform -1 0 3564 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_158
timestamp 1751266522
transform -1 0 3588 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_152
timestamp 1751266522
transform -1 0 3612 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_112
timestamp 1751266522
transform -1 0 3644 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_384
timestamp 1751266522
transform -1 0 3676 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_50
timestamp 1751266522
transform -1 0 3716 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_181
timestamp 1751266522
transform 1 0 3716 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_127
timestamp 1751266522
transform 1 0 3740 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_13
timestamp 1751266522
transform 1 0 3756 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_108
timestamp 1751266522
transform 1 0 3804 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_212
timestamp 1751266522
transform -1 0 3860 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_110
timestamp 1751266522
transform 1 0 3860 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_213
timestamp 1751266522
transform 1 0 3884 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1751266522
transform 1 0 3916 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_221
timestamp 1751266522
transform 1 0 3940 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_7_0
timestamp 1751266522
transform 1 0 3972 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_7_1
timestamp 1751266522
transform 1 0 3980 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_67
timestamp 1751266522
transform 1 0 3988 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_66
timestamp 1751266522
transform 1 0 4012 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_222
timestamp 1751266522
transform 1 0 4036 0 -1 2305
box -2 -3 34 103
use BUFX2  BUFX2_70
timestamp 1751266522
transform -1 0 4092 0 -1 2305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_3
timestamp 1751266522
transform -1 0 4148 0 -1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_194
timestamp 1751266522
transform -1 0 4180 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_55
timestamp 1751266522
transform 1 0 4180 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_49
timestamp 1751266522
transform -1 0 4220 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_183
timestamp 1751266522
transform -1 0 4252 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_91
timestamp 1751266522
transform 1 0 4252 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_98
timestamp 1751266522
transform -1 0 4292 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_60
timestamp 1751266522
transform -1 0 4316 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_181
timestamp 1751266522
transform 1 0 4316 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1751266522
transform -1 0 4380 0 -1 2305
box -2 -3 34 103
use FILL  FILL_23_1
timestamp 1751266522
transform -1 0 4388 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_2
timestamp 1751266522
transform -1 0 4396 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_16
timestamp 1751266522
transform -1 0 28 0 1 2305
box -2 -3 26 103
use DFFSR  DFFSR_64
timestamp 1751266522
transform -1 0 204 0 1 2305
box -2 -3 178 103
use CLKBUF1  CLKBUF1_13
timestamp 1751266522
transform 1 0 204 0 1 2305
box -2 -3 74 103
use DFFSR  DFFSR_58
timestamp 1751266522
transform 1 0 276 0 1 2305
box -2 -3 178 103
use FILL  FILL_23_0_0
timestamp 1751266522
transform 1 0 452 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1751266522
transform 1 0 460 0 1 2305
box -2 -3 10 103
use INVX1  INVX1_66
timestamp 1751266522
transform 1 0 468 0 1 2305
box -2 -3 18 103
use DFFSR  DFFSR_55
timestamp 1751266522
transform 1 0 484 0 1 2305
box -2 -3 178 103
use INVX2  INVX2_31
timestamp 1751266522
transform 1 0 660 0 1 2305
box -2 -3 18 103
use DFFSR  DFFSR_52
timestamp 1751266522
transform -1 0 852 0 1 2305
box -2 -3 178 103
use FILL  FILL_23_1_0
timestamp 1751266522
transform 1 0 852 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1751266522
transform 1 0 860 0 1 2305
box -2 -3 10 103
use DFFSR  DFFSR_53
timestamp 1751266522
transform 1 0 868 0 1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_98
timestamp 1751266522
transform 1 0 1044 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_54
timestamp 1751266522
transform -1 0 1108 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1751266522
transform -1 0 1140 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_33
timestamp 1751266522
transform -1 0 1156 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_41
timestamp 1751266522
transform 1 0 1156 0 1 2305
box -2 -3 34 103
use DFFSR  DFFSR_80
timestamp 1751266522
transform 1 0 1188 0 1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_67
timestamp 1751266522
transform -1 0 1396 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1751266522
transform 1 0 1396 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_2_0
timestamp 1751266522
transform 1 0 1420 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1751266522
transform 1 0 1428 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_5
timestamp 1751266522
transform 1 0 1436 0 1 2305
box -2 -3 26 103
use OAI22X1  OAI22X1_39
timestamp 1751266522
transform -1 0 1500 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_13
timestamp 1751266522
transform -1 0 1532 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1751266522
transform -1 0 1548 0 1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_12
timestamp 1751266522
transform 1 0 1548 0 1 2305
box -2 -3 74 103
use NOR2X1  NOR2X1_11
timestamp 1751266522
transform 1 0 1620 0 1 2305
box -2 -3 26 103
use OAI22X1  OAI22X1_28
timestamp 1751266522
transform 1 0 1644 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_46
timestamp 1751266522
transform -1 0 1700 0 1 2305
box -2 -3 18 103
use OAI22X1  OAI22X1_37
timestamp 1751266522
transform 1 0 1700 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_47
timestamp 1751266522
transform -1 0 1756 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_55
timestamp 1751266522
transform -1 0 1772 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_84
timestamp 1751266522
transform 1 0 1772 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_60
timestamp 1751266522
transform -1 0 1828 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_54
timestamp 1751266522
transform -1 0 1844 0 1 2305
box -2 -3 18 103
use AOI22X1  AOI22X1_25
timestamp 1751266522
transform 1 0 1844 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_174
timestamp 1751266522
transform 1 0 1884 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_3_0
timestamp 1751266522
transform 1 0 1916 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1751266522
transform 1 0 1924 0 1 2305
box -2 -3 10 103
use AOI22X1  AOI22X1_19
timestamp 1751266522
transform 1 0 1932 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_33
timestamp 1751266522
transform -1 0 2004 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1751266522
transform -1 0 2028 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_23
timestamp 1751266522
transform 1 0 2028 0 1 2305
box -2 -3 42 103
use OAI21X1  OAI21X1_321
timestamp 1751266522
transform -1 0 2100 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1751266522
transform 1 0 2100 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_320
timestamp 1751266522
transform 1 0 2132 0 1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_74
timestamp 1751266522
transform 1 0 2164 0 1 2305
box -2 -3 42 103
use NOR2X1  NOR2X1_127
timestamp 1751266522
transform -1 0 2228 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_126
timestamp 1751266522
transform -1 0 2252 0 1 2305
box -2 -3 26 103
use DFFSR  DFFSR_127
timestamp 1751266522
transform -1 0 2428 0 1 2305
box -2 -3 178 103
use FILL  FILL_23_4_0
timestamp 1751266522
transform 1 0 2428 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1751266522
transform 1 0 2436 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_637
timestamp 1751266522
transform 1 0 2444 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_238
timestamp 1751266522
transform 1 0 2476 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_641
timestamp 1751266522
transform -1 0 2532 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_220
timestamp 1751266522
transform 1 0 2532 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1751266522
transform -1 0 2588 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_236
timestamp 1751266522
transform 1 0 2588 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_92
timestamp 1751266522
transform 1 0 2612 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_635
timestamp 1751266522
transform 1 0 2628 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_591
timestamp 1751266522
transform -1 0 2692 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_58
timestamp 1751266522
transform 1 0 2692 0 1 2305
box -2 -3 18 103
use BUFX4  BUFX4_149
timestamp 1751266522
transform -1 0 2740 0 1 2305
box -2 -3 34 103
use INVX4  INVX4_10
timestamp 1751266522
transform -1 0 2764 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_475
timestamp 1751266522
transform 1 0 2764 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_59
timestamp 1751266522
transform 1 0 2796 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_423
timestamp 1751266522
transform 1 0 2812 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_476
timestamp 1751266522
transform 1 0 2844 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_424
timestamp 1751266522
transform 1 0 2876 0 1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_85
timestamp 1751266522
transform 1 0 2908 0 1 2305
box -2 -3 42 103
use FILL  FILL_23_5_0
timestamp 1751266522
transform -1 0 2956 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1751266522
transform -1 0 2964 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_139
timestamp 1751266522
transform -1 0 2996 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_422
timestamp 1751266522
transform -1 0 3028 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_167
timestamp 1751266522
transform 1 0 3028 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_361
timestamp 1751266522
transform -1 0 3084 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_5
timestamp 1751266522
transform 1 0 3084 0 1 2305
box -2 -3 50 103
use BUFX4  BUFX4_85
timestamp 1751266522
transform -1 0 3164 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_355
timestamp 1751266522
transform -1 0 3196 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_91
timestamp 1751266522
transform 1 0 3196 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_85
timestamp 1751266522
transform 1 0 3228 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_38
timestamp 1751266522
transform 1 0 3260 0 1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_84
timestamp 1751266522
transform 1 0 3300 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_354
timestamp 1751266522
transform -1 0 3364 0 1 2305
box -2 -3 34 103
use DFFSR  DFFSR_240
timestamp 1751266522
transform -1 0 3540 0 1 2305
box -2 -3 178 103
use FILL  FILL_23_6_0
timestamp 1751266522
transform -1 0 3548 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1751266522
transform -1 0 3556 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_385
timestamp 1751266522
transform -1 0 3588 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_113
timestamp 1751266522
transform 1 0 3588 0 1 2305
box -2 -3 34 103
use DFFSR  DFFSR_224
timestamp 1751266522
transform 1 0 3620 0 1 2305
box -2 -3 178 103
use NAND2X1  NAND2X1_109
timestamp 1751266522
transform 1 0 3796 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_101
timestamp 1751266522
transform 1 0 3820 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_59
timestamp 1751266522
transform -1 0 3868 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1751266522
transform 1 0 3868 0 1 2305
box -2 -3 26 103
use AND2X2  AND2X2_11
timestamp 1751266522
transform 1 0 3892 0 1 2305
box -2 -3 34 103
use XOR2X1  XOR2X1_6
timestamp 1751266522
transform 1 0 3924 0 1 2305
box -2 -3 58 103
use FILL  FILL_23_7_0
timestamp 1751266522
transform -1 0 3988 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_7_1
timestamp 1751266522
transform -1 0 3996 0 1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_73
timestamp 1751266522
transform -1 0 4020 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_182
timestamp 1751266522
transform -1 0 4052 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_129
timestamp 1751266522
transform -1 0 4076 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_132
timestamp 1751266522
transform 1 0 4076 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_131
timestamp 1751266522
transform -1 0 4124 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_196
timestamp 1751266522
transform 1 0 4124 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_85
timestamp 1751266522
transform 1 0 4156 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_195
timestamp 1751266522
transform 1 0 4172 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_252
timestamp 1751266522
transform 1 0 4204 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_128
timestamp 1751266522
transform -1 0 4260 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_80
timestamp 1751266522
transform 1 0 4260 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_95
timestamp 1751266522
transform -1 0 4308 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_180
timestamp 1751266522
transform 1 0 4308 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1751266522
transform -1 0 4364 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1751266522
transform 1 0 4364 0 1 2305
box -2 -3 34 103
use DFFSR  DFFSR_109
timestamp 1751266522
transform 1 0 4 0 -1 2505
box -2 -3 178 103
use NOR2X1  NOR2X1_21
timestamp 1751266522
transform 1 0 180 0 -1 2505
box -2 -3 26 103
use DFFSR  DFFSR_110
timestamp 1751266522
transform -1 0 380 0 -1 2505
box -2 -3 178 103
use INVX1  INVX1_75
timestamp 1751266522
transform 1 0 380 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_0_0
timestamp 1751266522
transform -1 0 404 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1751266522
transform -1 0 412 0 -1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_3
timestamp 1751266522
transform -1 0 484 0 -1 2505
box -2 -3 74 103
use INVX1  INVX1_73
timestamp 1751266522
transform -1 0 500 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_83
timestamp 1751266522
transform -1 0 524 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_184
timestamp 1751266522
transform -1 0 556 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1751266522
transform 1 0 556 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_31
timestamp 1751266522
transform 1 0 580 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_179
timestamp 1751266522
transform -1 0 636 0 -1 2505
box -2 -3 34 103
use DFFSR  DFFSR_50
timestamp 1751266522
transform -1 0 812 0 -1 2505
box -2 -3 178 103
use INVX2  INVX2_42
timestamp 1751266522
transform 1 0 812 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_1_0
timestamp 1751266522
transform 1 0 828 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1751266522
transform 1 0 836 0 -1 2505
box -2 -3 10 103
use DFFSR  DFFSR_59
timestamp 1751266522
transform 1 0 844 0 -1 2505
box -2 -3 178 103
use INVX2  INVX2_35
timestamp 1751266522
transform 1 0 1020 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_216
timestamp 1751266522
transform -1 0 1068 0 -1 2505
box -2 -3 34 103
use DFFSR  DFFSR_57
timestamp 1751266522
transform 1 0 1068 0 -1 2505
box -2 -3 178 103
use BUFX2  BUFX2_81
timestamp 1751266522
transform 1 0 1244 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1751266522
transform 1 0 1268 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1751266522
transform -1 0 1332 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1751266522
transform 1 0 1332 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_71
timestamp 1751266522
transform -1 0 1380 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_84
timestamp 1751266522
transform -1 0 1412 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_2_0
timestamp 1751266522
transform 1 0 1412 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1751266522
transform 1 0 1420 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_68
timestamp 1751266522
transform 1 0 1428 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_20
timestamp 1751266522
transform -1 0 1476 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_26
timestamp 1751266522
transform -1 0 1492 0 -1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_37
timestamp 1751266522
transform 1 0 1492 0 -1 2505
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1751266522
transform 1 0 1524 0 -1 2505
box -2 -3 42 103
use NAND3X1  NAND3X1_38
timestamp 1751266522
transform -1 0 1596 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_69
timestamp 1751266522
transform -1 0 1628 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1751266522
transform -1 0 1660 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1751266522
transform -1 0 1684 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_30
timestamp 1751266522
transform -1 0 1724 0 -1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_10
timestamp 1751266522
transform -1 0 1756 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_45
timestamp 1751266522
transform -1 0 1772 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_63
timestamp 1751266522
transform -1 0 1796 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_26
timestamp 1751266522
transform -1 0 1828 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1751266522
transform -1 0 1860 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_21
timestamp 1751266522
transform -1 0 1892 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1751266522
transform 1 0 1892 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_3_0
timestamp 1751266522
transform 1 0 1924 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1751266522
transform 1 0 1932 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_290
timestamp 1751266522
transform 1 0 1940 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_62
timestamp 1751266522
transform -1 0 2012 0 -1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_101
timestamp 1751266522
transform -1 0 2036 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_289
timestamp 1751266522
transform -1 0 2068 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_276
timestamp 1751266522
transform -1 0 2100 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_58
timestamp 1751266522
transform 1 0 2100 0 -1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_93
timestamp 1751266522
transform -1 0 2164 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_117
timestamp 1751266522
transform 1 0 2164 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_167
timestamp 1751266522
transform -1 0 2212 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_34
timestamp 1751266522
transform -1 0 2260 0 -1 2505
box -2 -3 50 103
use INVX1  INVX1_116
timestamp 1751266522
transform 1 0 2260 0 -1 2505
box -2 -3 18 103
use MUX2X1  MUX2X1_16
timestamp 1751266522
transform -1 0 2324 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_514
timestamp 1751266522
transform 1 0 2324 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1751266522
transform -1 0 2380 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_4_0
timestamp 1751266522
transform -1 0 2388 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1751266522
transform -1 0 2396 0 -1 2505
box -2 -3 10 103
use DFFSR  DFFSR_125
timestamp 1751266522
transform -1 0 2572 0 -1 2505
box -2 -3 178 103
use INVX1  INVX1_100
timestamp 1751266522
transform -1 0 2588 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_642
timestamp 1751266522
transform -1 0 2620 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_643
timestamp 1751266522
transform -1 0 2652 0 -1 2505
box -2 -3 34 103
use AND2X2  AND2X2_28
timestamp 1751266522
transform 1 0 2652 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_53
timestamp 1751266522
transform 1 0 2684 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_54
timestamp 1751266522
transform 1 0 2700 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_518
timestamp 1751266522
transform 1 0 2716 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_517
timestamp 1751266522
transform -1 0 2780 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_164
timestamp 1751266522
transform 1 0 2780 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_148
timestamp 1751266522
transform 1 0 2812 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_15
timestamp 1751266522
transform 1 0 2844 0 -1 2505
box -2 -3 50 103
use OAI22X1  OAI22X1_93
timestamp 1751266522
transform 1 0 2892 0 -1 2505
box -2 -3 42 103
use FILL  FILL_24_5_0
timestamp 1751266522
transform 1 0 2932 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1751266522
transform 1 0 2940 0 -1 2505
box -2 -3 10 103
use MUX2X1  MUX2X1_2
timestamp 1751266522
transform 1 0 2948 0 -1 2505
box -2 -3 50 103
use MUX2X1  MUX2X1_6
timestamp 1751266522
transform 1 0 2996 0 -1 2505
box -2 -3 50 103
use BUFX4  BUFX4_43
timestamp 1751266522
transform -1 0 3076 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_153
timestamp 1751266522
transform -1 0 3108 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_474
timestamp 1751266522
transform 1 0 3108 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_193
timestamp 1751266522
transform -1 0 3164 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_176
timestamp 1751266522
transform -1 0 3188 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_419
timestamp 1751266522
transform -1 0 3220 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_420
timestamp 1751266522
transform 1 0 3220 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_169
timestamp 1751266522
transform -1 0 3276 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_191
timestamp 1751266522
transform 1 0 3276 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_166
timestamp 1751266522
transform 1 0 3300 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_230
timestamp 1751266522
transform -1 0 3356 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_129
timestamp 1751266522
transform -1 0 3372 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_152
timestamp 1751266522
transform -1 0 3404 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1751266522
transform -1 0 3420 0 -1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_152
timestamp 1751266522
transform -1 0 3452 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_6_0
timestamp 1751266522
transform -1 0 3460 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1751266522
transform -1 0 3468 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_471
timestamp 1751266522
transform -1 0 3500 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_175
timestamp 1751266522
transform 1 0 3500 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_429
timestamp 1751266522
transform 1 0 3524 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_14
timestamp 1751266522
transform 1 0 3556 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_417
timestamp 1751266522
transform -1 0 3636 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_77
timestamp 1751266522
transform 1 0 3636 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_123
timestamp 1751266522
transform 1 0 3668 0 -1 2505
box -2 -3 34 103
use NOR3X1  NOR3X1_8
timestamp 1751266522
transform 1 0 3700 0 -1 2505
box -2 -3 66 103
use AOI21X1  AOI21X1_71
timestamp 1751266522
transform 1 0 3764 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_245
timestamp 1751266522
transform -1 0 3828 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_89
timestamp 1751266522
transform -1 0 3844 0 -1 2505
box -2 -3 18 103
use INVX4  INVX4_3
timestamp 1751266522
transform 1 0 3844 0 -1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_8
timestamp 1751266522
transform -1 0 3924 0 -1 2505
box -2 -3 58 103
use BUFX2  BUFX2_71
timestamp 1751266522
transform 1 0 3924 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_270
timestamp 1751266522
transform 1 0 3948 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_7_0
timestamp 1751266522
transform 1 0 3980 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_7_1
timestamp 1751266522
transform 1 0 3988 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_115
timestamp 1751266522
transform 1 0 3996 0 -1 2505
box -2 -3 26 103
use INVX8  INVX8_12
timestamp 1751266522
transform 1 0 4020 0 -1 2505
box -2 -3 42 103
use INVX4  INVX4_8
timestamp 1751266522
transform -1 0 4084 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_269
timestamp 1751266522
transform 1 0 4084 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_271
timestamp 1751266522
transform 1 0 4116 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_198
timestamp 1751266522
transform 1 0 4148 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_113
timestamp 1751266522
transform -1 0 4204 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_251
timestamp 1751266522
transform -1 0 4236 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_200
timestamp 1751266522
transform 1 0 4236 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_199
timestamp 1751266522
transform -1 0 4300 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_87
timestamp 1751266522
transform -1 0 4316 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_90
timestamp 1751266522
transform -1 0 4340 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1751266522
transform -1 0 4364 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_203
timestamp 1751266522
transform -1 0 4396 0 -1 2505
box -2 -3 34 103
use BUFX2  BUFX2_35
timestamp 1751266522
transform -1 0 28 0 1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_2
timestamp 1751266522
transform 1 0 28 0 1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_180
timestamp 1751266522
transform 1 0 84 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_47
timestamp 1751266522
transform -1 0 132 0 1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_23
timestamp 1751266522
transform 1 0 132 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1751266522
transform -1 0 180 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_181
timestamp 1751266522
transform 1 0 180 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1751266522
transform -1 0 236 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_182
timestamp 1751266522
transform -1 0 268 0 1 2505
box -2 -3 34 103
use DFFSR  DFFSR_111
timestamp 1751266522
transform -1 0 444 0 1 2505
box -2 -3 178 103
use FILL  FILL_25_0_0
timestamp 1751266522
transform -1 0 452 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1751266522
transform -1 0 460 0 1 2505
box -2 -3 10 103
use INVX8  INVX8_9
timestamp 1751266522
transform -1 0 500 0 1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_32
timestamp 1751266522
transform 1 0 500 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_89
timestamp 1751266522
transform -1 0 556 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_71
timestamp 1751266522
transform 1 0 556 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_35
timestamp 1751266522
transform 1 0 572 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_73
timestamp 1751266522
transform -1 0 620 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_34
timestamp 1751266522
transform -1 0 644 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1751266522
transform -1 0 660 0 1 2505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_22
timestamp 1751266522
transform -1 0 732 0 1 2505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_51
timestamp 1751266522
transform 1 0 732 0 1 2505
box -2 -3 74 103
use OAI21X1  OAI21X1_166
timestamp 1751266522
transform -1 0 836 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_164
timestamp 1751266522
transform -1 0 868 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_1_0
timestamp 1751266522
transform 1 0 868 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1751266522
transform 1 0 876 0 1 2505
box -2 -3 10 103
use DFFSR  DFFSR_63
timestamp 1751266522
transform 1 0 884 0 1 2505
box -2 -3 178 103
use INVX1  INVX1_64
timestamp 1751266522
transform 1 0 1060 0 1 2505
box -2 -3 18 103
use OAI22X1  OAI22X1_47
timestamp 1751266522
transform 1 0 1076 0 1 2505
box -2 -3 42 103
use INVX2  INVX2_22
timestamp 1751266522
transform -1 0 1132 0 1 2505
box -2 -3 18 103
use DFFSR  DFFSR_45
timestamp 1751266522
transform -1 0 1308 0 1 2505
box -2 -3 178 103
use DFFSR  DFFSR_36
timestamp 1751266522
transform 1 0 1308 0 1 2505
box -2 -3 178 103
use FILL  FILL_25_2_0
timestamp 1751266522
transform 1 0 1484 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1751266522
transform 1 0 1492 0 1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_20
timestamp 1751266522
transform 1 0 1500 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_36
timestamp 1751266522
transform -1 0 1556 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1751266522
transform -1 0 1588 0 1 2505
box -2 -3 34 103
use DFFSR  DFFSR_44
timestamp 1751266522
transform 1 0 1588 0 1 2505
box -2 -3 178 103
use INVX2  INVX2_18
timestamp 1751266522
transform -1 0 1780 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_21
timestamp 1751266522
transform 1 0 1780 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_18
timestamp 1751266522
transform 1 0 1804 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_20
timestamp 1751266522
transform 1 0 1828 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_92
timestamp 1751266522
transform -1 0 1892 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_25
timestamp 1751266522
transform 1 0 1892 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_3_0
timestamp 1751266522
transform 1 0 1924 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1751266522
transform 1 0 1932 0 1 2505
box -2 -3 10 103
use BUFX4  BUFX4_228
timestamp 1751266522
transform 1 0 1940 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_102
timestamp 1751266522
transform -1 0 1996 0 1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_21
timestamp 1751266522
transform -1 0 2044 0 1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_589
timestamp 1751266522
transform 1 0 2044 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_588
timestamp 1751266522
transform 1 0 2076 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_92
timestamp 1751266522
transform 1 0 2108 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_633
timestamp 1751266522
transform 1 0 2132 0 1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_22
timestamp 1751266522
transform -1 0 2212 0 1 2505
box -2 -3 50 103
use NOR2X1  NOR2X1_216
timestamp 1751266522
transform 1 0 2212 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_232
timestamp 1751266522
transform -1 0 2260 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_219
timestamp 1751266522
transform 1 0 2260 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_182
timestamp 1751266522
transform -1 0 2308 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_587
timestamp 1751266522
transform 1 0 2308 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_597
timestamp 1751266522
transform 1 0 2340 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_235
timestamp 1751266522
transform -1 0 2396 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_188
timestamp 1751266522
transform 1 0 2396 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_151
timestamp 1751266522
transform 1 0 2420 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_4_0
timestamp 1751266522
transform 1 0 2436 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1751266522
transform 1 0 2444 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_553
timestamp 1751266522
transform 1 0 2452 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_184
timestamp 1751266522
transform 1 0 2484 0 1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_105
timestamp 1751266522
transform 1 0 2508 0 1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_167
timestamp 1751266522
transform 1 0 2548 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_516
timestamp 1751266522
transform -1 0 2612 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_194
timestamp 1751266522
transform 1 0 2612 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_152
timestamp 1751266522
transform -1 0 2652 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_556
timestamp 1751266522
transform -1 0 2684 0 1 2505
box -2 -3 34 103
use DFFSR  DFFSR_191
timestamp 1751266522
transform -1 0 2860 0 1 2505
box -2 -3 178 103
use DFFSR  DFFSR_207
timestamp 1751266522
transform -1 0 3036 0 1 2505
box -2 -3 178 103
use FILL  FILL_25_5_0
timestamp 1751266522
transform 1 0 3036 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1751266522
transform 1 0 3044 0 1 2505
box -2 -3 10 103
use INVX2  INVX2_130
timestamp 1751266522
transform 1 0 3052 0 1 2505
box -2 -3 18 103
use BUFX4  BUFX4_44
timestamp 1751266522
transform 1 0 3068 0 1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_84
timestamp 1751266522
transform 1 0 3100 0 1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_196
timestamp 1751266522
transform -1 0 3164 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_138
timestamp 1751266522
transform -1 0 3196 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_418
timestamp 1751266522
transform -1 0 3228 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_178
timestamp 1751266522
transform -1 0 3252 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_472
timestamp 1751266522
transform -1 0 3284 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_473
timestamp 1751266522
transform 1 0 3284 0 1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_92
timestamp 1751266522
transform 1 0 3316 0 1 2505
box -2 -3 42 103
use DFFSR  DFFSR_192
timestamp 1751266522
transform -1 0 3532 0 1 2505
box -2 -3 178 103
use FILL  FILL_25_6_0
timestamp 1751266522
transform -1 0 3540 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1751266522
transform -1 0 3548 0 1 2505
box -2 -3 10 103
use NOR3X1  NOR3X1_9
timestamp 1751266522
transform -1 0 3612 0 1 2505
box -2 -3 66 103
use AOI21X1  AOI21X1_76
timestamp 1751266522
transform -1 0 3644 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_134
timestamp 1751266522
transform -1 0 3660 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_257
timestamp 1751266522
transform 1 0 3660 0 1 2505
box -2 -3 34 103
use AND2X2  AND2X2_13
timestamp 1751266522
transform -1 0 3724 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_9
timestamp 1751266522
transform -1 0 3756 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_247
timestamp 1751266522
transform 1 0 3756 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_125
timestamp 1751266522
transform -1 0 3812 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_57
timestamp 1751266522
transform -1 0 3836 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_69
timestamp 1751266522
transform 1 0 3836 0 1 2505
box -2 -3 26 103
use OR2X2  OR2X2_8
timestamp 1751266522
transform 1 0 3860 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_254
timestamp 1751266522
transform -1 0 3924 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_127
timestamp 1751266522
transform -1 0 3940 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_236
timestamp 1751266522
transform 1 0 3940 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_7_0
timestamp 1751266522
transform -1 0 3980 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_7_1
timestamp 1751266522
transform -1 0 3988 0 1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_63
timestamp 1751266522
transform -1 0 4020 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_257
timestamp 1751266522
transform 1 0 4020 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_130
timestamp 1751266522
transform 1 0 4052 0 1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_13
timestamp 1751266522
transform -1 0 4132 0 1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_234
timestamp 1751266522
transform 1 0 4132 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_235
timestamp 1751266522
transform -1 0 4196 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1751266522
transform -1 0 4220 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_61
timestamp 1751266522
transform 1 0 4220 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_72
timestamp 1751266522
transform 1 0 4244 0 1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_4
timestamp 1751266522
transform -1 0 4324 0 1 2505
box -2 -3 58 103
use BUFX2  BUFX2_73
timestamp 1751266522
transform -1 0 4348 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_91
timestamp 1751266522
transform -1 0 4372 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_96
timestamp 1751266522
transform -1 0 4396 0 1 2505
box -2 -3 26 103
use DFFSR  DFFSR_112
timestamp 1751266522
transform 1 0 4 0 -1 2705
box -2 -3 178 103
use NOR2X1  NOR2X1_46
timestamp 1751266522
transform 1 0 180 0 -1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_33
timestamp 1751266522
transform -1 0 244 0 -1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_185
timestamp 1751266522
transform -1 0 276 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1751266522
transform -1 0 300 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_22
timestamp 1751266522
transform -1 0 324 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_68
timestamp 1751266522
transform -1 0 348 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1751266522
transform 1 0 348 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1751266522
transform -1 0 396 0 -1 2705
box -2 -3 18 103
use FILL  FILL_26_0_0
timestamp 1751266522
transform -1 0 404 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1751266522
transform -1 0 412 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_47
timestamp 1751266522
transform -1 0 436 0 -1 2705
box -2 -3 26 103
use NOR3X1  NOR3X1_2
timestamp 1751266522
transform 1 0 436 0 -1 2705
box -2 -3 66 103
use OAI21X1  OAI21X1_183
timestamp 1751266522
transform 1 0 500 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_187
timestamp 1751266522
transform -1 0 564 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1751266522
transform -1 0 596 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_72
timestamp 1751266522
transform 1 0 596 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_33
timestamp 1751266522
transform 1 0 620 0 -1 2705
box -2 -3 26 103
use DFFSR  DFFSR_103
timestamp 1751266522
transform 1 0 644 0 -1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_167
timestamp 1751266522
transform -1 0 852 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_161
timestamp 1751266522
transform 1 0 852 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_68
timestamp 1751266522
transform 1 0 884 0 -1 2705
box -2 -3 18 103
use FILL  FILL_26_1_0
timestamp 1751266522
transform -1 0 908 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1751266522
transform -1 0 916 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_165
timestamp 1751266522
transform -1 0 948 0 -1 2705
box -2 -3 34 103
use DFFSR  DFFSR_102
timestamp 1751266522
transform -1 0 1124 0 -1 2705
box -2 -3 178 103
use BUFX2  BUFX2_69
timestamp 1751266522
transform 1 0 1124 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_212
timestamp 1751266522
transform 1 0 1148 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_90
timestamp 1751266522
transform -1 0 1212 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_76
timestamp 1751266522
transform -1 0 1244 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_33
timestamp 1751266522
transform -1 0 1268 0 -1 2705
box -2 -3 26 103
use DFFSR  DFFSR_43
timestamp 1751266522
transform 1 0 1268 0 -1 2705
box -2 -3 178 103
use FILL  FILL_26_2_0
timestamp 1751266522
transform 1 0 1444 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1751266522
transform 1 0 1452 0 -1 2705
box -2 -3 10 103
use DFFSR  DFFSR_66
timestamp 1751266522
transform 1 0 1460 0 -1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_66
timestamp 1751266522
transform -1 0 1668 0 -1 2705
box -2 -3 34 103
use DFFSR  DFFSR_42
timestamp 1751266522
transform 1 0 1668 0 -1 2705
box -2 -3 178 103
use BUFX4  BUFX4_23
timestamp 1751266522
transform -1 0 1876 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1751266522
transform 1 0 1876 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_88
timestamp 1751266522
transform 1 0 1908 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_3_0
timestamp 1751266522
transform -1 0 1948 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1751266522
transform -1 0 1956 0 -1 2705
box -2 -3 10 103
use DFFSR  DFFSR_144
timestamp 1751266522
transform -1 0 2132 0 -1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_634
timestamp 1751266522
transform 1 0 2132 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_33
timestamp 1751266522
transform -1 0 2212 0 -1 2705
box -2 -3 50 103
use NAND2X1  NAND2X1_225
timestamp 1751266522
transform -1 0 2236 0 -1 2705
box -2 -3 26 103
use OR2X2  OR2X2_10
timestamp 1751266522
transform -1 0 2268 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_132
timestamp 1751266522
transform 1 0 2268 0 -1 2705
box -2 -3 18 103
use OAI22X1  OAI22X1_104
timestamp 1751266522
transform 1 0 2284 0 -1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_515
timestamp 1751266522
transform -1 0 2356 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_513
timestamp 1751266522
transform -1 0 2388 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_166
timestamp 1751266522
transform -1 0 2420 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_192
timestamp 1751266522
transform 1 0 2420 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_4_0
timestamp 1751266522
transform 1 0 2444 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1751266522
transform 1 0 2452 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_554
timestamp 1751266522
transform 1 0 2460 0 -1 2705
box -2 -3 34 103
use DFFSR  DFFSR_159
timestamp 1751266522
transform -1 0 2668 0 -1 2705
box -2 -3 178 103
use NOR2X1  NOR2X1_209
timestamp 1751266522
transform -1 0 2692 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_557
timestamp 1751266522
transform 1 0 2692 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_114
timestamp 1751266522
transform -1 0 2764 0 -1 2705
box -2 -3 42 103
use INVX2  INVX2_79
timestamp 1751266522
transform 1 0 2764 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_561
timestamp 1751266522
transform 1 0 2780 0 -1 2705
box -2 -3 34 103
use DFFSR  DFFSR_208
timestamp 1751266522
transform -1 0 2988 0 -1 2705
box -2 -3 178 103
use FILL  FILL_26_5_0
timestamp 1751266522
transform 1 0 2988 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1751266522
transform 1 0 2996 0 -1 2705
box -2 -3 10 103
use INVX2  INVX2_82
timestamp 1751266522
transform 1 0 3004 0 -1 2705
box -2 -3 18 103
use INVX2  INVX2_81
timestamp 1751266522
transform 1 0 3020 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_431
timestamp 1751266522
transform 1 0 3036 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_87
timestamp 1751266522
transform 1 0 3068 0 -1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_432
timestamp 1751266522
transform -1 0 3140 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_481
timestamp 1751266522
transform -1 0 3172 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_141
timestamp 1751266522
transform 1 0 3172 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_430
timestamp 1751266522
transform -1 0 3236 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_155
timestamp 1751266522
transform 1 0 3236 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_480
timestamp 1751266522
transform 1 0 3268 0 -1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_7
timestamp 1751266522
transform -1 0 3348 0 -1 2705
box -2 -3 50 103
use DFFSR  DFFSR_247
timestamp 1751266522
transform 1 0 3348 0 -1 2705
box -2 -3 178 103
use FILL  FILL_26_6_0
timestamp 1751266522
transform 1 0 3524 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1751266522
transform 1 0 3532 0 -1 2705
box -2 -3 10 103
use OAI22X1  OAI22X1_121
timestamp 1751266522
transform 1 0 3540 0 -1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_703
timestamp 1751266522
transform -1 0 3612 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_255
timestamp 1751266522
transform 1 0 3612 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_272
timestamp 1751266522
transform -1 0 3668 0 -1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_34
timestamp 1751266522
transform 1 0 3668 0 -1 2705
box -2 -3 42 103
use NAND2X1  NAND2X1_135
timestamp 1751266522
transform 1 0 3708 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_256
timestamp 1751266522
transform -1 0 3764 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1751266522
transform -1 0 3788 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_121
timestamp 1751266522
transform 1 0 3788 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_255
timestamp 1751266522
transform 1 0 3812 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_84
timestamp 1751266522
transform -1 0 3860 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_54
timestamp 1751266522
transform 1 0 3860 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_253
timestamp 1751266522
transform 1 0 3884 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_122
timestamp 1751266522
transform 1 0 3916 0 -1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_265
timestamp 1751266522
transform -1 0 3972 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_7_0
timestamp 1751266522
transform -1 0 3980 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_7_1
timestamp 1751266522
transform -1 0 3988 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_68
timestamp 1751266522
transform -1 0 4020 0 -1 2705
box -2 -3 34 103
use INVX4  INVX4_4
timestamp 1751266522
transform -1 0 4044 0 -1 2705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_12
timestamp 1751266522
transform -1 0 4100 0 -1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_202
timestamp 1751266522
transform -1 0 4132 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_256
timestamp 1751266522
transform 1 0 4132 0 -1 2705
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1751266522
transform -1 0 4196 0 -1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_9
timestamp 1751266522
transform 1 0 4196 0 -1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_201
timestamp 1751266522
transform 1 0 4252 0 -1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1751266522
transform -1 0 4340 0 -1 2705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_5
timestamp 1751266522
transform -1 0 4396 0 -1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_188
timestamp 1751266522
transform -1 0 36 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1751266522
transform 1 0 36 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1751266522
transform 1 0 68 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1751266522
transform -1 0 124 0 1 2705
box -2 -3 26 103
use NOR3X1  NOR3X1_3
timestamp 1751266522
transform -1 0 188 0 1 2705
box -2 -3 66 103
use NAND2X1  NAND2X1_86
timestamp 1751266522
transform -1 0 212 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_78
timestamp 1751266522
transform -1 0 228 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_25
timestamp 1751266522
transform 1 0 228 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_77
timestamp 1751266522
transform -1 0 276 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_186
timestamp 1751266522
transform 1 0 276 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_0_0
timestamp 1751266522
transform -1 0 316 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1751266522
transform -1 0 324 0 1 2705
box -2 -3 10 103
use DFFSR  DFFSR_113
timestamp 1751266522
transform -1 0 500 0 1 2705
box -2 -3 178 103
use NAND2X1  NAND2X1_85
timestamp 1751266522
transform -1 0 524 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_160
timestamp 1751266522
transform 1 0 524 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_69
timestamp 1751266522
transform -1 0 572 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_178
timestamp 1751266522
transform 1 0 572 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_47
timestamp 1751266522
transform 1 0 604 0 1 2705
box -2 -3 74 103
use NAND2X1  NAND2X1_75
timestamp 1751266522
transform -1 0 700 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_38
timestamp 1751266522
transform 1 0 700 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_170
timestamp 1751266522
transform -1 0 756 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1751266522
transform -1 0 780 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_74
timestamp 1751266522
transform -1 0 804 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_5
timestamp 1751266522
transform -1 0 836 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_20
timestamp 1751266522
transform -1 0 868 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1751266522
transform 1 0 868 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_80
timestamp 1751266522
transform 1 0 892 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_1_0
timestamp 1751266522
transform -1 0 924 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1751266522
transform -1 0 932 0 1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_39
timestamp 1751266522
transform -1 0 956 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_6
timestamp 1751266522
transform -1 0 988 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_163
timestamp 1751266522
transform -1 0 1020 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1751266522
transform 1 0 1020 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_46
timestamp 1751266522
transform -1 0 1060 0 1 2705
box -2 -3 18 103
use DFFSR  DFFSR_54
timestamp 1751266522
transform -1 0 1236 0 1 2705
box -2 -3 178 103
use BUFX4  BUFX4_122
timestamp 1751266522
transform -1 0 1268 0 1 2705
box -2 -3 34 103
use DFFSR  DFFSR_41
timestamp 1751266522
transform 1 0 1268 0 1 2705
box -2 -3 178 103
use FILL  FILL_27_2_0
timestamp 1751266522
transform -1 0 1452 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1751266522
transform -1 0 1460 0 1 2705
box -2 -3 10 103
use BUFX2  BUFX2_51
timestamp 1751266522
transform -1 0 1484 0 1 2705
box -2 -3 26 103
use BUFX2  BUFX2_79
timestamp 1751266522
transform -1 0 1508 0 1 2705
box -2 -3 26 103
use DFFSR  DFFSR_74
timestamp 1751266522
transform -1 0 1684 0 1 2705
box -2 -3 178 103
use BUFX2  BUFX2_37
timestamp 1751266522
transform 1 0 1684 0 1 2705
box -2 -3 26 103
use DFFSR  DFFSR_93
timestamp 1751266522
transform -1 0 1884 0 1 2705
box -2 -3 178 103
use FILL  FILL_27_3_0
timestamp 1751266522
transform -1 0 1892 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1751266522
transform -1 0 1900 0 1 2705
box -2 -3 10 103
use DFFSR  DFFSR_176
timestamp 1751266522
transform -1 0 2076 0 1 2705
box -2 -3 178 103
use NAND3X1  NAND3X1_252
timestamp 1751266522
transform 1 0 2076 0 1 2705
box -2 -3 34 103
use MUX2X1  MUX2X1_25
timestamp 1751266522
transform 1 0 2108 0 1 2705
box -2 -3 50 103
use MUX2X1  MUX2X1_26
timestamp 1751266522
transform 1 0 2156 0 1 2705
box -2 -3 50 103
use OAI21X1  OAI21X1_598
timestamp 1751266522
transform -1 0 2236 0 1 2705
box -2 -3 34 103
use DFFSR  DFFSR_141
timestamp 1751266522
transform 1 0 2236 0 1 2705
box -2 -3 178 103
use INVX2  INVX2_131
timestamp 1751266522
transform 1 0 2412 0 1 2705
box -2 -3 18 103
use FILL  FILL_27_4_0
timestamp 1751266522
transform 1 0 2428 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1751266522
transform 1 0 2436 0 1 2705
box -2 -3 10 103
use OAI22X1  OAI22X1_113
timestamp 1751266522
transform 1 0 2444 0 1 2705
box -2 -3 42 103
use INVX4  INVX4_9
timestamp 1751266522
transform 1 0 2484 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_208
timestamp 1751266522
transform -1 0 2532 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_185
timestamp 1751266522
transform 1 0 2532 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_552
timestamp 1751266522
transform 1 0 2564 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_197
timestamp 1751266522
transform 1 0 2596 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_153
timestamp 1751266522
transform 1 0 2620 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_522
timestamp 1751266522
transform -1 0 2668 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_210
timestamp 1751266522
transform -1 0 2692 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_186
timestamp 1751266522
transform 1 0 2692 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_555
timestamp 1751266522
transform 1 0 2724 0 1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_115
timestamp 1751266522
transform 1 0 2756 0 1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_562
timestamp 1751266522
transform -1 0 2828 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_189
timestamp 1751266522
transform 1 0 2828 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_560
timestamp 1751266522
transform -1 0 2892 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1751266522
transform -1 0 2900 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1751266522
transform -1 0 2908 0 1 2705
box -2 -3 10 103
use DFFSR  DFFSR_189
timestamp 1751266522
transform -1 0 3084 0 1 2705
box -2 -3 178 103
use OAI22X1  OAI22X1_95
timestamp 1751266522
transform 1 0 3084 0 1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_482
timestamp 1751266522
transform -1 0 3156 0 1 2705
box -2 -3 34 103
use DFFSR  DFFSR_246
timestamp 1751266522
transform 1 0 3156 0 1 2705
box -2 -3 178 103
use XNOR2X1  XNOR2X1_14
timestamp 1751266522
transform 1 0 3332 0 1 2705
box -2 -3 58 103
use AOI21X1  AOI21X1_222
timestamp 1751266522
transform 1 0 3388 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_254
timestamp 1751266522
transform 1 0 3420 0 1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_276
timestamp 1751266522
transform -1 0 3476 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_6_0
timestamp 1751266522
transform 1 0 3476 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1751266522
transform 1 0 3484 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_707
timestamp 1751266522
transform 1 0 3492 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_260
timestamp 1751266522
transform 1 0 3524 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_50
timestamp 1751266522
transform 1 0 3548 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_60
timestamp 1751266522
transform 1 0 3564 0 1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_6
timestamp 1751266522
transform -1 0 3652 0 1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_248
timestamp 1751266522
transform 1 0 3652 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_127
timestamp 1751266522
transform 1 0 3684 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_70
timestamp 1751266522
transform -1 0 3740 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_76
timestamp 1751266522
transform -1 0 3764 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_128
timestamp 1751266522
transform -1 0 3780 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_94
timestamp 1751266522
transform -1 0 3804 0 1 2705
box -2 -3 26 103
use OR2X2  OR2X2_4
timestamp 1751266522
transform -1 0 3836 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_209
timestamp 1751266522
transform -1 0 3868 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_48
timestamp 1751266522
transform -1 0 3892 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1751266522
transform 1 0 3892 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_242
timestamp 1751266522
transform 1 0 3924 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_67
timestamp 1751266522
transform 1 0 3956 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_7_0
timestamp 1751266522
transform 1 0 3988 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_7_1
timestamp 1751266522
transform 1 0 3996 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_197
timestamp 1751266522
transform 1 0 4004 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1751266522
transform 1 0 4036 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_87
timestamp 1751266522
transform -1 0 4084 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_9
timestamp 1751266522
transform -1 0 4116 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_88
timestamp 1751266522
transform -1 0 4132 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_88
timestamp 1751266522
transform -1 0 4156 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_10
timestamp 1751266522
transform 1 0 4156 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_253
timestamp 1751266522
transform -1 0 4220 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_211
timestamp 1751266522
transform -1 0 4252 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_49
timestamp 1751266522
transform -1 0 4276 0 1 2705
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1751266522
transform -1 0 4300 0 1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_222
timestamp 1751266522
transform 1 0 4300 0 1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_4
timestamp 1751266522
transform -1 0 4388 0 1 2705
box -2 -3 58 103
use FILL  FILL_28_1
timestamp 1751266522
transform 1 0 4388 0 1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_23
timestamp 1751266522
transform -1 0 28 0 -1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_5
timestamp 1751266522
transform 1 0 28 0 -1 2905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_67
timestamp 1751266522
transform 1 0 100 0 -1 2905
box -2 -3 74 103
use INVX1  INVX1_80
timestamp 1751266522
transform 1 0 172 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_189
timestamp 1751266522
transform 1 0 188 0 -1 2905
box -2 -3 34 103
use OAI22X1  OAI22X1_50
timestamp 1751266522
transform -1 0 260 0 -1 2905
box -2 -3 42 103
use INVX1  INVX1_79
timestamp 1751266522
transform -1 0 276 0 -1 2905
box -2 -3 18 103
use DFFSR  DFFSR_100
timestamp 1751266522
transform 1 0 276 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_0_0
timestamp 1751266522
transform 1 0 452 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1751266522
transform 1 0 460 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_158
timestamp 1751266522
transform 1 0 468 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_77
timestamp 1751266522
transform -1 0 524 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_90
timestamp 1751266522
transform -1 0 556 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_72
timestamp 1751266522
transform 1 0 556 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_177
timestamp 1751266522
transform -1 0 604 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1751266522
transform 1 0 604 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1751266522
transform -1 0 660 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_108
timestamp 1751266522
transform -1 0 836 0 -1 2905
box -2 -3 178 103
use NAND2X1  NAND2X1_78
timestamp 1751266522
transform -1 0 860 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_88
timestamp 1751266522
transform 1 0 860 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_65
timestamp 1751266522
transform -1 0 908 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_1_0
timestamp 1751266522
transform -1 0 916 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1751266522
transform -1 0 924 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_162
timestamp 1751266522
transform -1 0 956 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_173
timestamp 1751266522
transform 1 0 956 0 -1 2905
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1751266522
transform 1 0 988 0 -1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_175
timestamp 1751266522
transform -1 0 1076 0 -1 2905
box -2 -3 34 103
use INVX8  INVX8_10
timestamp 1751266522
transform 1 0 1076 0 -1 2905
box -2 -3 42 103
use CLKBUF1  CLKBUF1_39
timestamp 1751266522
transform -1 0 1188 0 -1 2905
box -2 -3 74 103
use DFFSR  DFFSR_39
timestamp 1751266522
transform 1 0 1188 0 -1 2905
box -2 -3 178 103
use INVX2  INVX2_29
timestamp 1751266522
transform 1 0 1364 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_76
timestamp 1751266522
transform 1 0 1380 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_2_0
timestamp 1751266522
transform -1 0 1412 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1751266522
transform -1 0 1420 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_19
timestamp 1751266522
transform -1 0 1452 0 -1 2905
box -2 -3 34 103
use BUFX2  BUFX2_77
timestamp 1751266522
transform -1 0 1476 0 -1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_26
timestamp 1751266522
transform -1 0 1548 0 -1 2905
box -2 -3 74 103
use BUFX2  BUFX2_45
timestamp 1751266522
transform 1 0 1548 0 -1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_18
timestamp 1751266522
transform -1 0 1644 0 -1 2905
box -2 -3 74 103
use NAND3X1  NAND3X1_42
timestamp 1751266522
transform -1 0 1676 0 -1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_30
timestamp 1751266522
transform -1 0 1748 0 -1 2905
box -2 -3 74 103
use BUFX4  BUFX4_119
timestamp 1751266522
transform 1 0 1748 0 -1 2905
box -2 -3 34 103
use MUX2X1  MUX2X1_1
timestamp 1751266522
transform 1 0 1780 0 -1 2905
box -2 -3 50 103
use NOR2X1  NOR2X1_52
timestamp 1751266522
transform 1 0 1828 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_3_0
timestamp 1751266522
transform 1 0 1852 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1751266522
transform 1 0 1860 0 -1 2905
box -2 -3 10 103
use DFFSR  DFFSR_65
timestamp 1751266522
transform 1 0 1868 0 -1 2905
box -2 -3 178 103
use INVX1  INVX1_82
timestamp 1751266522
transform 1 0 2044 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_232
timestamp 1751266522
transform 1 0 2060 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_128
timestamp 1751266522
transform 1 0 2092 0 -1 2905
box -2 -3 178 103
use OAI21X1  OAI21X1_281
timestamp 1751266522
transform -1 0 2300 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_136
timestamp 1751266522
transform -1 0 2316 0 -1 2905
box -2 -3 18 103
use INVX2  INVX2_80
timestamp 1751266522
transform 1 0 2316 0 -1 2905
box -2 -3 18 103
use DFFSR  DFFSR_160
timestamp 1751266522
transform -1 0 2508 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_4_0
timestamp 1751266522
transform 1 0 2508 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1751266522
transform 1 0 2516 0 -1 2905
box -2 -3 10 103
use OAI22X1  OAI22X1_106
timestamp 1751266522
transform 1 0 2524 0 -1 2905
box -2 -3 42 103
use AOI21X1  AOI21X1_170
timestamp 1751266522
transform -1 0 2596 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_521
timestamp 1751266522
transform 1 0 2596 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_523
timestamp 1751266522
transform -1 0 2660 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_157
timestamp 1751266522
transform -1 0 2836 0 -1 2905
box -2 -3 178 103
use NOR2X1  NOR2X1_51
timestamp 1751266522
transform 1 0 2836 0 -1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_29
timestamp 1751266522
transform 1 0 2860 0 -1 2905
box -2 -3 74 103
use NOR2X1  NOR2X1_258
timestamp 1751266522
transform 1 0 2932 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_5_0
timestamp 1751266522
transform -1 0 2964 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1751266522
transform -1 0 2972 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_81
timestamp 1751266522
transform -1 0 2988 0 -1 2905
box -2 -3 18 103
use DFFSR  DFFSR_205
timestamp 1751266522
transform -1 0 3164 0 -1 2905
box -2 -3 178 103
use NAND2X1  NAND2X1_259
timestamp 1751266522
transform 1 0 3164 0 -1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_90
timestamp 1751266522
transform -1 0 3228 0 -1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_710
timestamp 1751266522
transform -1 0 3260 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1751266522
transform -1 0 3284 0 -1 2905
box -2 -3 26 103
use DFFSR  DFFSR_251
timestamp 1751266522
transform 1 0 3284 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_6_0
timestamp 1751266522
transform 1 0 3460 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1751266522
transform 1 0 3468 0 -1 2905
box -2 -3 10 103
use OAI22X1  OAI22X1_122
timestamp 1751266522
transform 1 0 3476 0 -1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_704
timestamp 1751266522
transform -1 0 3548 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_256
timestamp 1751266522
transform 1 0 3548 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_258
timestamp 1751266522
transform 1 0 3572 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_709
timestamp 1751266522
transform 1 0 3596 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1751266522
transform 1 0 3628 0 -1 2905
box -2 -3 26 103
use OAI22X1  OAI22X1_123
timestamp 1751266522
transform -1 0 3692 0 -1 2905
box -2 -3 42 103
use INVX2  INVX2_51
timestamp 1751266522
transform 1 0 3692 0 -1 2905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_10
timestamp 1751266522
transform -1 0 3764 0 -1 2905
box -2 -3 58 103
use INVX1  INVX1_126
timestamp 1751266522
transform 1 0 3764 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_240
timestamp 1751266522
transform -1 0 3812 0 -1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_6
timestamp 1751266522
transform -1 0 3876 0 -1 2905
box -2 -3 66 103
use NAND3X1  NAND3X1_262
timestamp 1751266522
transform 1 0 3876 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1751266522
transform -1 0 3940 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_250
timestamp 1751266522
transform -1 0 3972 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_7_0
timestamp 1751266522
transform -1 0 3980 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_7_1
timestamp 1751266522
transform -1 0 3988 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_75
timestamp 1751266522
transform -1 0 4020 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_131
timestamp 1751266522
transform -1 0 4036 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_261
timestamp 1751266522
transform 1 0 4036 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_126
timestamp 1751266522
transform 1 0 4068 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_249
timestamp 1751266522
transform -1 0 4124 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1751266522
transform 1 0 4124 0 -1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_11
timestamp 1751266522
transform -1 0 4204 0 -1 2905
box -2 -3 58 103
use INVX2  INVX2_52
timestamp 1751266522
transform 1 0 4204 0 -1 2905
box -2 -3 18 103
use NOR3X1  NOR3X1_5
timestamp 1751266522
transform 1 0 4220 0 -1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_204
timestamp 1751266522
transform 1 0 4284 0 -1 2905
box -2 -3 34 103
use INVX4  INVX4_6
timestamp 1751266522
transform 1 0 4316 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_205
timestamp 1751266522
transform 1 0 4340 0 -1 2905
box -2 -3 34 103
use FILL  FILL_29_1
timestamp 1751266522
transform -1 0 4380 0 -1 2905
box -2 -3 10 103
use FILL  FILL_29_2
timestamp 1751266522
transform -1 0 4388 0 -1 2905
box -2 -3 10 103
use FILL  FILL_29_3
timestamp 1751266522
transform -1 0 4396 0 -1 2905
box -2 -3 10 103
use DFFSR  DFFSR_114
timestamp 1751266522
transform -1 0 180 0 1 2905
box -2 -3 178 103
use DFFSR  DFFSR_115
timestamp 1751266522
transform 1 0 180 0 1 2905
box -2 -3 178 103
use NAND2X1  NAND2X1_69
timestamp 1751266522
transform 1 0 356 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1751266522
transform -1 0 404 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_0_0
timestamp 1751266522
transform 1 0 404 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1751266522
transform 1 0 412 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_25
timestamp 1751266522
transform 1 0 420 0 1 2905
box -2 -3 26 103
use OR2X2  OR2X2_2
timestamp 1751266522
transform 1 0 444 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_235
timestamp 1751266522
transform 1 0 476 0 1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1751266522
transform -1 0 572 0 1 2905
box -2 -3 66 103
use AND2X2  AND2X2_4
timestamp 1751266522
transform -1 0 604 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1751266522
transform 1 0 604 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1751266522
transform 1 0 628 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_40
timestamp 1751266522
transform 1 0 652 0 1 2905
box -2 -3 26 103
use DFFSR  DFFSR_107
timestamp 1751266522
transform -1 0 852 0 1 2905
box -2 -3 178 103
use NOR2X1  NOR2X1_29
timestamp 1751266522
transform 1 0 852 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1751266522
transform 1 0 876 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_1_0
timestamp 1751266522
transform 1 0 908 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1751266522
transform 1 0 916 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_176
timestamp 1751266522
transform 1 0 924 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1751266522
transform 1 0 956 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_71
timestamp 1751266522
transform 1 0 980 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_238
timestamp 1751266522
transform -1 0 1036 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_101
timestamp 1751266522
transform -1 0 1212 0 1 2905
box -2 -3 178 103
use DFFSR  DFFSR_97
timestamp 1751266522
transform 1 0 1212 0 1 2905
box -2 -3 178 103
use OAI22X1  OAI22X1_48
timestamp 1751266522
transform -1 0 1428 0 1 2905
box -2 -3 42 103
use FILL  FILL_29_2_0
timestamp 1751266522
transform 1 0 1428 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1751266522
transform 1 0 1436 0 1 2905
box -2 -3 10 103
use OAI22X1  OAI22X1_49
timestamp 1751266522
transform 1 0 1444 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_190
timestamp 1751266522
transform 1 0 1484 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_191
timestamp 1751266522
transform -1 0 1548 0 1 2905
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1751266522
transform 1 0 1548 0 1 2905
box -2 -3 34 103
use OR2X2  OR2X2_3
timestamp 1751266522
transform -1 0 1612 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_98
timestamp 1751266522
transform 1 0 1612 0 1 2905
box -2 -3 178 103
use DFFSR  DFFSR_76
timestamp 1751266522
transform -1 0 1964 0 1 2905
box -2 -3 178 103
use FILL  FILL_29_3_0
timestamp 1751266522
transform 1 0 1964 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1751266522
transform 1 0 1972 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_44
timestamp 1751266522
transform 1 0 1980 0 1 2905
box -2 -3 74 103
use BUFX2  BUFX2_36
timestamp 1751266522
transform 1 0 2052 0 1 2905
box -2 -3 26 103
use DFFSR  DFFSR_244
timestamp 1751266522
transform -1 0 2252 0 1 2905
box -2 -3 178 103
use NAND2X1  NAND2X1_139
timestamp 1751266522
transform 1 0 2252 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_280
timestamp 1751266522
transform -1 0 2308 0 1 2905
box -2 -3 34 103
use BUFX2  BUFX2_76
timestamp 1751266522
transform -1 0 2332 0 1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_48
timestamp 1751266522
transform -1 0 2404 0 1 2905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_49
timestamp 1751266522
transform -1 0 2476 0 1 2905
box -2 -3 74 103
use FILL  FILL_29_4_0
timestamp 1751266522
transform 1 0 2476 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1751266522
transform 1 0 2484 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_2
timestamp 1751266522
transform 1 0 2492 0 1 2905
box -2 -3 74 103
use NOR2X1  NOR2X1_263
timestamp 1751266522
transform -1 0 2588 0 1 2905
box -2 -3 26 103
use DFFSR  DFFSR_245
timestamp 1751266522
transform 1 0 2588 0 1 2905
box -2 -3 178 103
use AOI21X1  AOI21X1_224
timestamp 1751266522
transform -1 0 2796 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_262
timestamp 1751266522
transform -1 0 2820 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_262
timestamp 1751266522
transform -1 0 2844 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_711
timestamp 1751266522
transform 1 0 2844 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_223
timestamp 1751266522
transform 1 0 2876 0 1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_28
timestamp 1751266522
transform 1 0 2908 0 1 2905
box -2 -3 74 103
use FILL  FILL_29_5_0
timestamp 1751266522
transform 1 0 2980 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1751266522
transform 1 0 2988 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_33
timestamp 1751266522
transform 1 0 2996 0 1 2905
box -2 -3 74 103
use BUFX4  BUFX4_15
timestamp 1751266522
transform 1 0 3068 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_259
timestamp 1751266522
transform -1 0 3124 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_261
timestamp 1751266522
transform 1 0 3124 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_708
timestamp 1751266522
transform -1 0 3180 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_706
timestamp 1751266522
transform -1 0 3212 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_252
timestamp 1751266522
transform 1 0 3212 0 1 2905
box -2 -3 178 103
use INVX1  INVX1_158
timestamp 1751266522
transform 1 0 3388 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_261
timestamp 1751266522
transform 1 0 3404 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_275
timestamp 1751266522
transform 1 0 3428 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_6_0
timestamp 1751266522
transform -1 0 3468 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1751266522
transform -1 0 3476 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_260
timestamp 1751266522
transform -1 0 3500 0 1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_3
timestamp 1751266522
transform -1 0 3556 0 1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_705
timestamp 1751266522
transform 1 0 3556 0 1 2905
box -2 -3 34 103
use BUFX2  BUFX2_78
timestamp 1751266522
transform 1 0 3588 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_73
timestamp 1751266522
transform 1 0 3612 0 1 2905
box -2 -3 34 103
use BUFX2  BUFX2_74
timestamp 1751266522
transform -1 0 3668 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_74
timestamp 1751266522
transform 1 0 3668 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_271
timestamp 1751266522
transform 1 0 3700 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_266
timestamp 1751266522
transform 1 0 3732 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_65
timestamp 1751266522
transform -1 0 3796 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_125
timestamp 1751266522
transform -1 0 3812 0 1 2905
box -2 -3 18 103
use NOR3X1  NOR3X1_7
timestamp 1751266522
transform -1 0 3876 0 1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_241
timestamp 1751266522
transform 1 0 3876 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_66
timestamp 1751266522
transform -1 0 3940 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_117
timestamp 1751266522
transform -1 0 3964 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_7_0
timestamp 1751266522
transform -1 0 3972 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_7_1
timestamp 1751266522
transform -1 0 3980 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_243
timestamp 1751266522
transform -1 0 4012 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1751266522
transform -1 0 4036 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_62
timestamp 1751266522
transform -1 0 4068 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1751266522
transform -1 0 4100 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_255
timestamp 1751266522
transform 1 0 4100 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_258
timestamp 1751266522
transform -1 0 4164 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_263
timestamp 1751266522
transform -1 0 4196 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_116
timestamp 1751266522
transform 1 0 4196 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_118
timestamp 1751266522
transform -1 0 4244 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_124
timestamp 1751266522
transform -1 0 4260 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_233
timestamp 1751266522
transform -1 0 4292 0 1 2905
box -2 -3 34 103
use OR2X2  OR2X2_7
timestamp 1751266522
transform -1 0 4324 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_237
timestamp 1751266522
transform 1 0 4324 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_260
timestamp 1751266522
transform 1 0 4356 0 1 2905
box -2 -3 34 103
use FILL  FILL_30_1
timestamp 1751266522
transform 1 0 4388 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_55
timestamp 1751266522
transform 1 0 4 0 -1 3105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_34
timestamp 1751266522
transform 1 0 76 0 -1 3105
box -2 -3 74 103
use DFFSR  DFFSR_105
timestamp 1751266522
transform 1 0 148 0 -1 3105
box -2 -3 178 103
use BUFX4  BUFX4_237
timestamp 1751266522
transform -1 0 356 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_0_0
timestamp 1751266522
transform 1 0 356 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1751266522
transform 1 0 364 0 -1 3105
box -2 -3 10 103
use DFFSR  DFFSR_104
timestamp 1751266522
transform 1 0 372 0 -1 3105
box -2 -3 178 103
use OAI21X1  OAI21X1_169
timestamp 1751266522
transform 1 0 548 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_168
timestamp 1751266522
transform -1 0 612 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_42
timestamp 1751266522
transform -1 0 636 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_70
timestamp 1751266522
transform 1 0 636 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_41
timestamp 1751266522
transform 1 0 652 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_82
timestamp 1751266522
transform 1 0 676 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_171
timestamp 1751266522
transform 1 0 700 0 -1 3105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_1
timestamp 1751266522
transform -1 0 788 0 -1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_81
timestamp 1751266522
transform -1 0 812 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_27
timestamp 1751266522
transform 1 0 812 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_172
timestamp 1751266522
transform 1 0 836 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1751266522
transform 1 0 868 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_1_0
timestamp 1751266522
transform 1 0 900 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_1
timestamp 1751266522
transform 1 0 908 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_174
timestamp 1751266522
transform 1 0 916 0 -1 3105
box -2 -3 34 103
use DFFSR  DFFSR_106
timestamp 1751266522
transform -1 0 1124 0 -1 3105
box -2 -3 178 103
use BUFX4  BUFX4_236
timestamp 1751266522
transform -1 0 1156 0 -1 3105
box -2 -3 34 103
use INVX8  INVX8_11
timestamp 1751266522
transform -1 0 1196 0 -1 3105
box -2 -3 42 103
use INVX8  INVX8_8
timestamp 1751266522
transform 1 0 1196 0 -1 3105
box -2 -3 42 103
use INVX8  INVX8_26
timestamp 1751266522
transform -1 0 1276 0 -1 3105
box -2 -3 42 103
use DFFSR  DFFSR_99
timestamp 1751266522
transform 1 0 1276 0 -1 3105
box -2 -3 178 103
use FILL  FILL_30_2_0
timestamp 1751266522
transform -1 0 1460 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_1
timestamp 1751266522
transform -1 0 1468 0 -1 3105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_64
timestamp 1751266522
transform -1 0 1540 0 -1 3105
box -2 -3 74 103
use DFFSR  DFFSR_68
timestamp 1751266522
transform 1 0 1540 0 -1 3105
box -2 -3 178 103
use BUFX2  BUFX2_39
timestamp 1751266522
transform 1 0 1716 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_64
timestamp 1751266522
transform 1 0 1740 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_47
timestamp 1751266522
transform -1 0 1788 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1751266522
transform 1 0 1788 0 -1 3105
box -2 -3 26 103
use DFFSR  DFFSR_70
timestamp 1751266522
transform 1 0 1812 0 -1 3105
box -2 -3 178 103
use FILL  FILL_30_3_0
timestamp 1751266522
transform 1 0 1988 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_1
timestamp 1751266522
transform 1 0 1996 0 -1 3105
box -2 -3 10 103
use BUFX2  BUFX2_41
timestamp 1751266522
transform 1 0 2004 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1751266522
transform 1 0 2028 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_14
timestamp 1751266522
transform 1 0 2052 0 -1 3105
box -2 -3 34 103
use DFFSR  DFFSR_173
timestamp 1751266522
transform -1 0 2260 0 -1 3105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_37
timestamp 1751266522
transform -1 0 2332 0 -1 3105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_56
timestamp 1751266522
transform -1 0 2404 0 -1 3105
box -2 -3 74 103
use FILL  FILL_30_4_0
timestamp 1751266522
transform -1 0 2412 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_1
timestamp 1751266522
transform -1 0 2420 0 -1 3105
box -2 -3 10 103
use DFFSR  DFFSR_175
timestamp 1751266522
transform -1 0 2596 0 -1 3105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_41
timestamp 1751266522
transform -1 0 2668 0 -1 3105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_61
timestamp 1751266522
transform 1 0 2668 0 -1 3105
box -2 -3 74 103
use DFFSR  DFFSR_253
timestamp 1751266522
transform -1 0 2916 0 -1 3105
box -2 -3 178 103
use FILL  FILL_30_5_0
timestamp 1751266522
transform 1 0 2916 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_1
timestamp 1751266522
transform 1 0 2924 0 -1 3105
box -2 -3 10 103
use DFFSR  DFFSR_249
timestamp 1751266522
transform 1 0 2932 0 -1 3105
box -2 -3 178 103
use DFFSR  DFFSR_250
timestamp 1751266522
transform 1 0 3108 0 -1 3105
box -2 -3 178 103
use DFFSR  DFFSR_248
timestamp 1751266522
transform 1 0 3284 0 -1 3105
box -2 -3 178 103
use FILL  FILL_30_6_0
timestamp 1751266522
transform -1 0 3468 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_6_1
timestamp 1751266522
transform -1 0 3476 0 -1 3105
box -2 -3 10 103
use NAND3X1  NAND3X1_269
timestamp 1751266522
transform -1 0 3508 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_272
timestamp 1751266522
transform -1 0 3540 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_129
timestamp 1751266522
transform -1 0 3556 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_273
timestamp 1751266522
transform -1 0 3588 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_260
timestamp 1751266522
transform -1 0 3620 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_246
timestamp 1751266522
transform -1 0 3652 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_151
timestamp 1751266522
transform 1 0 3652 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_124
timestamp 1751266522
transform -1 0 3692 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_69
timestamp 1751266522
transform 1 0 3692 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1751266522
transform -1 0 3756 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_267
timestamp 1751266522
transform 1 0 3756 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1751266522
transform -1 0 3812 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_268
timestamp 1751266522
transform 1 0 3812 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1751266522
transform -1 0 3876 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_270
timestamp 1751266522
transform -1 0 3908 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1751266522
transform 1 0 3908 0 -1 3105
box -2 -3 26 103
use AND2X2  AND2X2_12
timestamp 1751266522
transform -1 0 3964 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1751266522
transform 1 0 3964 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_7_0
timestamp 1751266522
transform -1 0 3996 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_7_1
timestamp 1751266522
transform -1 0 4004 0 -1 3105
box -2 -3 10 103
use NAND3X1  NAND3X1_264
timestamp 1751266522
transform -1 0 4036 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_48
timestamp 1751266522
transform 1 0 4036 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_239
timestamp 1751266522
transform -1 0 4084 0 -1 3105
box -2 -3 34 103
use INVX4  INVX4_7
timestamp 1751266522
transform -1 0 4108 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_254
timestamp 1751266522
transform 1 0 4108 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_238
timestamp 1751266522
transform 1 0 4140 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_259
timestamp 1751266522
transform 1 0 4172 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_210
timestamp 1751266522
transform -1 0 4236 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1751266522
transform 1 0 4236 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_52
timestamp 1751266522
transform 1 0 4268 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_121
timestamp 1751266522
transform 1 0 4300 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_136
timestamp 1751266522
transform -1 0 4364 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_1
timestamp 1751266522
transform -1 0 4372 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_2
timestamp 1751266522
transform -1 0 4380 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_3
timestamp 1751266522
transform -1 0 4388 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_4
timestamp 1751266522
transform -1 0 4396 0 -1 3105
box -2 -3 10 103
<< labels >>
flabel metal6 s 392 -30 408 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 896 -30 912 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 138 -22 142 7 FreeSans 24 0 0 0 wb_clk_i
port 2 nsew
flabel metal2 s 1254 3128 1258 3132 3 FreeSans 24 90 0 0 wb_rst_i
port 3 nsew
flabel metal2 s 3694 -22 3698 -18 7 FreeSans 24 270 0 0 wb_adr_i[0]
port 4 nsew
flabel metal2 s 1638 3128 1642 3132 3 FreeSans 24 90 0 0 wb_adr_i[1]
port 5 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 wb_adr_i[2]
port 6 nsew
flabel metal3 s -26 1528 -22 1532 7 FreeSans 24 0 0 0 wb_adr_i[3]
port 7 nsew
flabel metal3 s -26 1488 -22 1492 7 FreeSans 24 0 0 0 wb_adr_i[4]
port 8 nsew
flabel metal2 s 2566 -22 2570 -18 7 FreeSans 24 270 0 0 wb_dat_i[0]
port 9 nsew
flabel metal3 s -26 1788 -22 1792 7 FreeSans 24 0 0 0 wb_dat_i[1]
port 10 nsew
flabel metal2 s 1438 -22 1442 -18 7 FreeSans 24 270 0 0 wb_dat_i[2]
port 11 nsew
flabel metal2 s 2750 -22 2754 -18 7 FreeSans 24 270 0 0 wb_dat_i[3]
port 12 nsew
flabel metal2 s 2638 -22 2642 -18 7 FreeSans 24 270 0 0 wb_dat_i[4]
port 13 nsew
flabel metal3 s -26 1648 -22 1652 7 FreeSans 24 0 0 0 wb_dat_i[5]
port 14 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 wb_dat_i[6]
port 15 nsew
flabel metal3 s -26 1178 -22 1182 7 FreeSans 24 0 0 0 wb_dat_i[7]
port 16 nsew
flabel metal2 s 1158 3128 1162 3132 3 FreeSans 24 90 0 0 wb_dat_i[8]
port 17 nsew
flabel metal2 s 2406 3128 2410 3132 3 FreeSans 24 90 0 0 wb_dat_i[9]
port 18 nsew
flabel metal2 s 1358 3128 1362 3132 3 FreeSans 24 90 0 0 wb_dat_i[10]
port 19 nsew
flabel metal2 s 2486 3128 2490 3132 3 FreeSans 24 90 0 0 wb_dat_i[11]
port 20 nsew
flabel metal2 s 2174 3128 2178 3132 3 FreeSans 24 90 0 0 wb_dat_i[12]
port 21 nsew
flabel metal2 s 2638 3128 2642 3132 3 FreeSans 24 90 0 0 wb_dat_i[13]
port 22 nsew
flabel metal3 s -26 1468 -22 1472 7 FreeSans 24 0 0 0 wb_dat_i[14]
port 23 nsew
flabel metal3 s -26 1448 -22 1452 7 FreeSans 24 0 0 0 wb_dat_i[15]
port 24 nsew
flabel metal2 s 2022 -22 2026 -18 7 FreeSans 24 270 0 0 wb_dat_i[16]
port 25 nsew
flabel metal2 s 2134 -22 2138 -18 7 FreeSans 24 270 0 0 wb_dat_i[17]
port 26 nsew
flabel metal2 s 2166 -22 2170 -18 7 FreeSans 24 270 0 0 wb_dat_i[18]
port 27 nsew
flabel metal2 s 2294 -22 2298 -18 7 FreeSans 24 270 0 0 wb_dat_i[19]
port 28 nsew
flabel metal2 s 2310 -22 2314 -18 7 FreeSans 24 270 0 0 wb_dat_i[20]
port 29 nsew
flabel metal2 s 1598 -22 1602 -18 7 FreeSans 24 270 0 0 wb_dat_i[21]
port 30 nsew
flabel metal2 s 1198 -22 1202 -18 7 FreeSans 24 270 0 0 wb_dat_i[22]
port 31 nsew
flabel metal2 s 2398 -22 2402 -18 7 FreeSans 24 270 0 0 wb_dat_i[23]
port 32 nsew
flabel metal3 s -26 1298 -22 1302 7 FreeSans 24 0 0 0 wb_dat_i[24]
port 33 nsew
flabel metal2 s 2142 3128 2146 3132 3 FreeSans 24 90 0 0 wb_dat_i[25]
port 34 nsew
flabel metal2 s 1006 -22 1010 -18 7 FreeSans 24 270 0 0 wb_dat_i[26]
port 35 nsew
flabel metal2 s 2566 3128 2570 3132 3 FreeSans 24 90 0 0 wb_dat_i[27]
port 36 nsew
flabel metal2 s 1998 3128 2002 3132 3 FreeSans 24 90 0 0 wb_dat_i[28]
port 37 nsew
flabel metal3 s -26 1278 -22 1282 7 FreeSans 24 0 0 0 wb_dat_i[29]
port 38 nsew
flabel metal2 s 2150 -22 2154 -18 7 FreeSans 24 270 0 0 wb_dat_i[30]
port 39 nsew
flabel metal2 s 1374 -22 1378 -18 7 FreeSans 24 270 0 0 wb_dat_i[31]
port 40 nsew
flabel metal3 s -26 748 -22 752 7 FreeSans 24 0 0 0 wb_sel_i[0]
port 41 nsew
flabel metal2 s 1902 3128 1906 3132 3 FreeSans 24 90 0 0 wb_sel_i[1]
port 42 nsew
flabel metal2 s 2270 -22 2274 -18 7 FreeSans 24 270 0 0 wb_sel_i[2]
port 43 nsew
flabel metal2 s 1918 3128 1922 3132 3 FreeSans 24 90 0 0 wb_sel_i[3]
port 44 nsew
flabel metal3 s -26 2268 -22 2272 7 FreeSans 24 0 0 0 wb_we_i
port 45 nsew
flabel metal3 s -26 2308 -22 2312 7 FreeSans 24 0 0 0 wb_stb_i
port 46 nsew
flabel metal3 s -26 2248 -22 2252 7 FreeSans 24 0 0 0 wb_cyc_i
port 47 nsew
flabel metal2 s 2246 3128 2250 3132 3 FreeSans 24 90 0 0 miso_pad_i
port 48 nsew
flabel metal2 s 2062 3128 2066 3132 3 FreeSans 24 90 0 0 wb_dat_o[0]
port 49 nsew
flabel metal2 s 1694 3128 1698 3132 3 FreeSans 24 90 0 0 wb_dat_o[1]
port 50 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 wb_dat_o[2]
port 51 nsew
flabel metal2 s 1726 3128 1730 3132 3 FreeSans 24 90 0 0 wb_dat_o[3]
port 52 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 wb_dat_o[4]
port 53 nsew
flabel metal2 s 2014 3128 2018 3132 3 FreeSans 24 90 0 0 wb_dat_o[5]
port 54 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 wb_dat_o[6]
port 55 nsew
flabel metal3 s -26 988 -22 992 7 FreeSans 24 0 0 0 wb_dat_o[7]
port 56 nsew
flabel metal2 s 558 -22 562 -18 7 FreeSans 24 270 0 0 wb_dat_o[8]
port 57 nsew
flabel metal2 s 1558 3128 1562 3132 3 FreeSans 24 90 0 0 wb_dat_o[9]
port 58 nsew
flabel metal3 s -26 1688 -22 1692 7 FreeSans 24 0 0 0 wb_dat_o[10]
port 59 nsew
flabel metal2 s 1774 3128 1778 3132 3 FreeSans 24 90 0 0 wb_dat_o[11]
port 60 nsew
flabel metal3 s -26 2288 -22 2292 7 FreeSans 24 0 0 0 wb_dat_o[12]
port 61 nsew
flabel metal3 s -26 1868 -22 1872 7 FreeSans 24 0 0 0 wb_dat_o[13]
port 62 nsew
flabel metal3 s -26 1388 -22 1392 7 FreeSans 24 0 0 0 wb_dat_o[14]
port 63 nsew
flabel metal2 s 1470 3128 1474 3132 3 FreeSans 24 90 0 0 wb_dat_o[15]
port 64 nsew
flabel metal3 s -26 68 -22 72 7 FreeSans 24 0 0 0 wb_dat_o[16]
port 65 nsew
flabel metal2 s 574 -22 578 -18 7 FreeSans 24 270 0 0 wb_dat_o[17]
port 66 nsew
flabel metal2 s 414 -22 418 -18 7 FreeSans 24 270 0 0 wb_dat_o[18]
port 67 nsew
flabel metal3 s -26 788 -22 792 7 FreeSans 24 0 0 0 wb_dat_o[19]
port 68 nsew
flabel metal2 s 358 -22 362 -18 7 FreeSans 24 270 0 0 wb_dat_o[20]
port 69 nsew
flabel metal2 s 1358 -22 1362 -18 7 FreeSans 24 270 0 0 wb_dat_o[21]
port 70 nsew
flabel metal3 s -26 348 -22 352 7 FreeSans 24 0 0 0 wb_dat_o[22]
port 71 nsew
flabel metal2 s 446 -22 450 -18 7 FreeSans 24 270 0 0 wb_dat_o[23]
port 72 nsew
flabel metal2 s 238 -22 242 -18 7 FreeSans 24 270 0 0 wb_dat_o[24]
port 73 nsew
flabel metal3 s -26 2148 -22 2152 7 FreeSans 24 0 0 0 wb_dat_o[25]
port 74 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 wb_dat_o[26]
port 75 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 wb_dat_o[27]
port 76 nsew
flabel metal2 s 1750 3128 1754 3132 3 FreeSans 24 90 0 0 wb_dat_o[28]
port 77 nsew
flabel metal3 s -26 1768 -22 1772 7 FreeSans 24 0 0 0 wb_dat_o[29]
port 78 nsew
flabel metal2 s 790 -22 794 -18 7 FreeSans 24 270 0 0 wb_dat_o[30]
port 79 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 wb_dat_o[31]
port 80 nsew
flabel metal3 s -26 2548 -22 2552 7 FreeSans 24 0 0 0 wb_ack_o
port 81 nsew
flabel metal2 s 4054 -22 4058 -18 7 FreeSans 24 270 0 0 wb_err_o
port 82 nsew
flabel metal2 s 1134 3128 1138 3132 3 FreeSans 24 90 0 0 wb_int_o
port 83 nsew
flabel metal3 s -26 1748 -22 1752 7 FreeSans 24 0 0 0 ss_pad_o[0]
port 84 nsew
flabel metal3 s -26 2048 -22 2052 7 FreeSans 24 0 0 0 ss_pad_o[1]
port 85 nsew
flabel metal3 s -26 848 -22 852 7 FreeSans 24 0 0 0 ss_pad_o[2]
port 86 nsew
flabel metal3 s -26 1968 -22 1972 7 FreeSans 24 0 0 0 ss_pad_o[3]
port 87 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 ss_pad_o[4]
port 88 nsew
flabel metal3 s -26 2008 -22 2012 7 FreeSans 24 0 0 0 ss_pad_o[5]
port 89 nsew
flabel metal3 s -26 1848 -22 1852 7 FreeSans 24 0 0 0 ss_pad_o[6]
port 90 nsew
flabel metal3 s -26 1508 -22 1512 7 FreeSans 24 0 0 0 ss_pad_o[7]
port 91 nsew
flabel metal3 s -26 1368 -22 1372 7 FreeSans 24 0 0 0 ss_pad_o[8]
port 92 nsew
flabel metal3 s -26 1068 -22 1072 7 FreeSans 24 0 0 0 ss_pad_o[9]
port 93 nsew
flabel metal3 s -26 1948 -22 1952 7 FreeSans 24 0 0 0 ss_pad_o[10]
port 94 nsew
flabel metal2 s 430 -22 434 -18 7 FreeSans 24 270 0 0 ss_pad_o[11]
port 95 nsew
flabel metal3 s -26 2188 -22 2192 7 FreeSans 24 0 0 0 ss_pad_o[12]
port 96 nsew
flabel metal3 s -26 1588 -22 1592 7 FreeSans 24 0 0 0 ss_pad_o[13]
port 97 nsew
flabel metal3 s -26 968 -22 972 7 FreeSans 24 0 0 0 ss_pad_o[14]
port 98 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 0 0 0 ss_pad_o[15]
port 99 nsew
flabel metal2 s 958 -22 962 -18 7 FreeSans 24 270 0 0 ss_pad_o[16]
port 100 nsew
flabel metal2 s 1070 -22 1074 -18 7 FreeSans 24 270 0 0 ss_pad_o[17]
port 101 nsew
flabel metal2 s 982 -22 986 -18 7 FreeSans 24 270 0 0 ss_pad_o[18]
port 102 nsew
flabel metal2 s 374 -22 378 -18 7 FreeSans 24 270 0 0 ss_pad_o[19]
port 103 nsew
flabel metal2 s 774 -22 778 -18 7 FreeSans 24 270 0 0 ss_pad_o[20]
port 104 nsew
flabel metal2 s 326 -22 330 -18 7 FreeSans 24 270 0 0 ss_pad_o[21]
port 105 nsew
flabel metal2 s 886 -22 890 -18 7 FreeSans 24 270 0 0 ss_pad_o[22]
port 106 nsew
flabel metal2 s 654 -22 658 -18 7 FreeSans 24 270 0 0 ss_pad_o[23]
port 107 nsew
flabel metal3 s -26 768 -22 772 7 FreeSans 24 0 0 0 ss_pad_o[24]
port 108 nsew
flabel metal3 s -26 1988 -22 1992 7 FreeSans 24 0 0 0 ss_pad_o[25]
port 109 nsew
flabel metal2 s 342 -22 346 -18 7 FreeSans 24 270 0 0 ss_pad_o[26]
port 110 nsew
flabel metal3 s -26 1668 -22 1672 7 FreeSans 24 0 0 0 ss_pad_o[27]
port 111 nsew
flabel metal3 s -26 2168 -22 2172 7 FreeSans 24 0 0 0 ss_pad_o[28]
port 112 nsew
flabel metal3 s -26 1568 -22 1572 7 FreeSans 24 0 0 0 ss_pad_o[29]
port 113 nsew
flabel metal2 s 542 -22 546 -18 7 FreeSans 24 270 0 0 ss_pad_o[30]
port 114 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 ss_pad_o[31]
port 115 nsew
flabel metal2 s 1798 3128 1802 3132 3 FreeSans 24 90 0 0 sclk_pad_o
port 116 nsew
flabel metal2 s 2038 3128 2042 3132 3 FreeSans 24 90 0 0 mosi_pad_o
port 117 nsew
<< end >>
