module spi_top ( gnd, vdd, wb_clk_i, wb_rst_i, wb_adr_i, wb_dat_i, wb_sel_i, wb_we_i, wb_stb_i, wb_cyc_i, miso_pad_i, wb_dat_o, wb_ack_o, wb_err_o, wb_int_o, ss_pad_o, sclk_pad_o, mosi_pad_o);

input gnd, vdd;
input wb_clk_i;
input wb_rst_i;
input wb_we_i;
input wb_stb_i;
input wb_cyc_i;
input miso_pad_i;
output wb_ack_o;
output wb_err_o;
output wb_int_o;
output sclk_pad_o;
output mosi_pad_o;
input [4:0] wb_adr_i;
input [31:0] wb_dat_i;
input [3:0] wb_sel_i;
output [31:0] wb_dat_o;
output [31:0] ss_pad_o;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf10), .Y(wb_clk_i_bF_buf10_bF_buf3) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf10), .Y(wb_clk_i_bF_buf10_bF_buf2) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf10), .Y(wb_clk_i_bF_buf10_bF_buf1) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf10), .Y(wb_clk_i_bF_buf10_bF_buf0) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf11), .Y(wb_clk_i_bF_buf11_bF_buf3) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf11), .Y(wb_clk_i_bF_buf11_bF_buf2) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf11), .Y(wb_clk_i_bF_buf11_bF_buf1) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf11), .Y(wb_clk_i_bF_buf11_bF_buf0) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf12), .Y(wb_clk_i_bF_buf12_bF_buf3) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf12), .Y(wb_clk_i_bF_buf12_bF_buf2) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf12), .Y(wb_clk_i_bF_buf12_bF_buf1) );
CLKBUF1 CLKBUF1_12 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf12), .Y(wb_clk_i_bF_buf12_bF_buf0) );
CLKBUF1 CLKBUF1_13 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf13), .Y(wb_clk_i_bF_buf13_bF_buf3) );
CLKBUF1 CLKBUF1_14 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf13), .Y(wb_clk_i_bF_buf13_bF_buf2) );
CLKBUF1 CLKBUF1_15 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf13), .Y(wb_clk_i_bF_buf13_bF_buf1) );
CLKBUF1 CLKBUF1_16 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf13), .Y(wb_clk_i_bF_buf13_bF_buf0) );
CLKBUF1 CLKBUF1_17 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf14), .Y(wb_clk_i_bF_buf14_bF_buf3) );
CLKBUF1 CLKBUF1_18 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf14), .Y(wb_clk_i_bF_buf14_bF_buf2) );
CLKBUF1 CLKBUF1_19 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf14), .Y(wb_clk_i_bF_buf14_bF_buf1) );
CLKBUF1 CLKBUF1_20 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf14), .Y(wb_clk_i_bF_buf14_bF_buf0) );
CLKBUF1 CLKBUF1_21 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf2), .Y(wb_clk_i_bF_buf2_bF_buf3) );
CLKBUF1 CLKBUF1_22 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf2), .Y(wb_clk_i_bF_buf2_bF_buf2) );
CLKBUF1 CLKBUF1_23 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf2), .Y(wb_clk_i_bF_buf2_bF_buf1) );
CLKBUF1 CLKBUF1_24 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf2), .Y(wb_clk_i_bF_buf2_bF_buf0) );
CLKBUF1 CLKBUF1_25 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf3), .Y(wb_clk_i_bF_buf3_bF_buf3) );
CLKBUF1 CLKBUF1_26 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf3), .Y(wb_clk_i_bF_buf3_bF_buf2) );
CLKBUF1 CLKBUF1_27 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf3), .Y(wb_clk_i_bF_buf3_bF_buf1) );
CLKBUF1 CLKBUF1_28 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf3), .Y(wb_clk_i_bF_buf3_bF_buf0) );
CLKBUF1 CLKBUF1_29 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf4), .Y(wb_clk_i_bF_buf4_bF_buf3) );
CLKBUF1 CLKBUF1_30 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf4), .Y(wb_clk_i_bF_buf4_bF_buf2) );
CLKBUF1 CLKBUF1_31 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf4), .Y(wb_clk_i_bF_buf4_bF_buf1) );
CLKBUF1 CLKBUF1_32 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf4), .Y(wb_clk_i_bF_buf4_bF_buf0) );
CLKBUF1 CLKBUF1_33 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf5), .Y(wb_clk_i_bF_buf5_bF_buf3) );
CLKBUF1 CLKBUF1_34 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf5), .Y(wb_clk_i_bF_buf5_bF_buf2) );
CLKBUF1 CLKBUF1_35 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf5), .Y(wb_clk_i_bF_buf5_bF_buf1) );
CLKBUF1 CLKBUF1_36 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf5), .Y(wb_clk_i_bF_buf5_bF_buf0) );
CLKBUF1 CLKBUF1_37 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf6), .Y(wb_clk_i_bF_buf6_bF_buf3) );
CLKBUF1 CLKBUF1_38 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf6), .Y(wb_clk_i_bF_buf6_bF_buf2) );
CLKBUF1 CLKBUF1_39 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf6), .Y(wb_clk_i_bF_buf6_bF_buf1) );
CLKBUF1 CLKBUF1_40 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf6), .Y(wb_clk_i_bF_buf6_bF_buf0) );
CLKBUF1 CLKBUF1_41 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf7), .Y(wb_clk_i_bF_buf7_bF_buf3) );
CLKBUF1 CLKBUF1_42 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf7), .Y(wb_clk_i_bF_buf7_bF_buf2) );
CLKBUF1 CLKBUF1_43 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf7), .Y(wb_clk_i_bF_buf7_bF_buf1) );
CLKBUF1 CLKBUF1_44 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf7), .Y(wb_clk_i_bF_buf7_bF_buf0) );
CLKBUF1 CLKBUF1_45 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf8), .Y(wb_clk_i_bF_buf8_bF_buf3) );
CLKBUF1 CLKBUF1_46 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf8), .Y(wb_clk_i_bF_buf8_bF_buf2) );
CLKBUF1 CLKBUF1_47 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf8), .Y(wb_clk_i_bF_buf8_bF_buf1) );
CLKBUF1 CLKBUF1_48 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf8), .Y(wb_clk_i_bF_buf8_bF_buf0) );
CLKBUF1 CLKBUF1_49 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf9), .Y(wb_clk_i_bF_buf9_bF_buf3) );
CLKBUF1 CLKBUF1_50 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf9), .Y(wb_clk_i_bF_buf9_bF_buf2) );
CLKBUF1 CLKBUF1_51 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf9), .Y(wb_clk_i_bF_buf9_bF_buf1) );
CLKBUF1 CLKBUF1_52 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i_bF_buf9), .Y(wb_clk_i_bF_buf9_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf6) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf5) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf4) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf3) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf2) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf1) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .Y(_1066__bF_buf0) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf10) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf9) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf8) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf7) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf6) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf5) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf4) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf3) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf2) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf1) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_547_), .Y(_547__bF_buf0) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf7_) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf6_) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf5_) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf4_) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf3_) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf2_) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf1_) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[1]), .Y(wb_sel_i_1_bF_buf0_) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf4) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf3) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf2) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf1) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf0) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .Y(_2094__bF_buf3) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .Y(_2094__bF_buf2) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .Y(_2094__bF_buf1) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .Y(_2094__bF_buf0) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .Y(_2091__bF_buf3) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .Y(_2091__bF_buf2) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .Y(_2091__bF_buf1) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .Y(_2091__bF_buf0) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf5) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf4) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf3) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf2) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf1) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_693__bF_buf0) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf5) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf4) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf3) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf2) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf1) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1606__bF_buf0) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_687_), .Y(_687__bF_buf3) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_687_), .Y(_687__bF_buf2) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_687_), .Y(_687__bF_buf1) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_687_), .Y(_687__bF_buf0) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf5) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf4) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf3) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf2) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf1) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .Y(_1603__bF_buf0) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1582__bF_buf4) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1582__bF_buf3) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1582__bF_buf2) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1582__bF_buf1) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .Y(_1582__bF_buf0) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_358_), .Y(_358__bF_buf3) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_358_), .Y(_358__bF_buf2) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_358_), .Y(_358__bF_buf1) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_358_), .Y(_358__bF_buf0) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf5) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf4) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf3) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf2) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf1) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1600__bF_buf0) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .Y(_2041__bF_buf3) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .Y(_2041__bF_buf2) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .Y(_2041__bF_buf1) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .Y(_2041__bF_buf0) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .Y(_1576__bF_buf4) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .Y(_1576__bF_buf3) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .Y(_1576__bF_buf2) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .Y(_1576__bF_buf1) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .Y(_1576__bF_buf0) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf6_) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf5_) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf4_) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf3_) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf2_) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf1_) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[3]), .Y(wb_sel_i_3_bF_buf0_) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf6) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf5) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf4) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf3) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf2) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf1) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_9__bF_buf0) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_12__bF_buf4) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_12__bF_buf3) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_12__bF_buf2) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_12__bF_buf1) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_12__bF_buf0) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf7_) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf6_) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf5_) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf4_) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf3_) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf2_) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf1_) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[0]), .Y(wb_sel_i_0_bF_buf0_) );
CLKBUF1 CLKBUF1_53 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf14) );
CLKBUF1 CLKBUF1_54 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf13) );
CLKBUF1 CLKBUF1_55 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf12) );
CLKBUF1 CLKBUF1_56 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf11) );
CLKBUF1 CLKBUF1_57 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf10) );
CLKBUF1 CLKBUF1_58 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf9) );
CLKBUF1 CLKBUF1_59 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf8) );
CLKBUF1 CLKBUF1_60 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf7) );
CLKBUF1 CLKBUF1_61 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf6) );
CLKBUF1 CLKBUF1_62 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf5) );
CLKBUF1 CLKBUF1_63 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf4) );
CLKBUF1 CLKBUF1_64 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf3) );
CLKBUF1 CLKBUF1_65 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf2) );
CLKBUF1 CLKBUF1_66 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf1) );
CLKBUF1 CLKBUF1_67 ( .gnd(gnd), .vdd(vdd), .A(wb_clk_i), .Y(wb_clk_i_bF_buf0) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_249__bF_buf4) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_249__bF_buf3) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_249__bF_buf2) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_249__bF_buf1) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_249__bF_buf0) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf9) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf8) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf7) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf6) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf5) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf4) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf3) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf2) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf1) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable), .Y(clgen_enable_bF_buf0) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_190__bF_buf3) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_190__bF_buf2) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_190__bF_buf1) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_190__bF_buf0) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf3) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf2) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf1) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_243__bF_buf0) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf6) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf5) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf4) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf3) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf2) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf1) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1561__bF_buf0) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_789__bF_buf3) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_789__bF_buf2) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_789__bF_buf1) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_789__bF_buf0) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1073__bF_buf4) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1073__bF_buf3) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1073__bF_buf2) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1073__bF_buf1) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1073__bF_buf0) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf8) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf7) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf6) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf5) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf4) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf3) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf2) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf1) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_686_), .Y(_686__bF_buf0) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf6) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf5) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf4) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf3) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf2) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf1) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .Y(_1067__bF_buf0) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .Y(_2081__bF_buf3) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .Y(_2081__bF_buf2) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .Y(_2081__bF_buf1) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .Y(_2081__bF_buf0) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf7) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf6) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf5) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf4) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf3) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf2) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf1) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2078__bF_buf0) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .Y(_1502__bF_buf3) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .Y(_1502__bF_buf2) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .Y(_1502__bF_buf1) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .Y(_1502__bF_buf0) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf6_) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf5_) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf4_) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf3_) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf2_) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf1_) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i[2]), .Y(wb_sel_i_2_bF_buf0_) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf3) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf2) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf1) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf0) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf7) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf6) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf5) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf4) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf3) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf2) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf1) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_11__bF_buf0) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1569__bF_buf4) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1569__bF_buf3) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1569__bF_buf2) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1569__bF_buf1) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1569__bF_buf0) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf8) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf7) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf6) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf5) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf4) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf3) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf2) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf1) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_5__bF_buf0) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_189__bF_buf3) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_189__bF_buf2) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_189__bF_buf1) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_189__bF_buf0) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf7) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf6) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf5) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf4) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf3) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf2) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf1) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .Y(_2025__bF_buf0) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf5) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf4) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf3) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf2) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf1) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf0) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(_433_), .Y(_433__bF_buf3) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(_433_), .Y(_433__bF_buf2) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(_433_), .Y(_433__bF_buf1) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(_433_), .Y(_433__bF_buf0) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(_242__bF_buf3) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(_242__bF_buf2) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(_242__bF_buf1) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(_242__bF_buf0) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf7) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf6) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf5) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf4) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf3) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf2) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf1) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_694__bF_buf0) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_788__bF_buf4) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_788__bF_buf3) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_788__bF_buf2) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_788__bF_buf1) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_788_), .Y(_788__bF_buf0) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .Y(_1072__bF_buf4) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .Y(_1072__bF_buf3) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .Y(_1072__bF_buf2) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .Y(_1072__bF_buf1) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .Y(_1072__bF_buf0) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf7) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf6) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf5) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf4) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf3) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf2) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf1) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_688_), .Y(_688__bF_buf0) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(lsb), .Y(lsb_bF_buf3) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(lsb), .Y(lsb_bF_buf2) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(lsb), .Y(lsb_bF_buf1) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(lsb), .Y(lsb_bF_buf0) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_685__bF_buf4) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_685__bF_buf3) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_685__bF_buf2) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_685__bF_buf1) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_685__bF_buf0) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(ss_24_), .Y(_6_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[2]), .Y(_7_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[4]), .B(wb_adr_i[3]), .C(_7_), .Y(_8_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf3), .Y(_9_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(wb_we_i), .B(wb_stb_i), .C(wb_cyc_i), .Y(_10_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_10_), .Y(_11_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf6), .B(_11__bF_buf7), .Y(_12_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[24]), .B(wb_sel_i_3_bF_buf6_), .Y(_13_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(wb_sel_i_3_bF_buf5_), .C(_13_), .Y(_14_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_14_), .C(_9__bF_buf5), .Y(_15_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_6_), .C(_15_), .Y(_2__24_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(ss_25_), .Y(_16_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf4_), .B(wb_dat_i[25]), .Y(_17_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(wb_sel_i_3_bF_buf3_), .C(_17_), .Y(_18_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_18_), .C(_9__bF_buf4), .Y(_19_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_16_), .C(_19_), .Y(_2__25_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(ss_26_), .Y(_20_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf2_), .B(wb_dat_i[26]), .Y(_21_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(wb_sel_i_3_bF_buf1_), .C(_21_), .Y(_22_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_22_), .C(_9__bF_buf3), .Y(_23_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_20_), .C(_23_), .Y(_2__26_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(ss_27_), .Y(_24_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf0_), .B(wb_dat_i[27]), .Y(_25_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(wb_sel_i_3_bF_buf6_), .C(_25_), .Y(_26_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_26_), .C(_9__bF_buf2), .Y(_27_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_24_), .C(_27_), .Y(_2__27_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(ss_28_), .Y(_28_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf5_), .B(wb_dat_i[28]), .Y(_29_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(wb_sel_i_3_bF_buf4_), .C(_29_), .Y(_30_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_30_), .C(_9__bF_buf1), .Y(_31_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_28_), .C(_31_), .Y(_2__28_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(ss_29_), .Y(_32_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf3_), .B(wb_dat_i[29]), .Y(_33_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(wb_sel_i_3_bF_buf2_), .C(_33_), .Y(_34_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_34_), .C(_9__bF_buf0), .Y(_35_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_32_), .C(_35_), .Y(_2__29_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(ss_30_), .Y(_36_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf1_), .B(wb_dat_i[30]), .Y(_37_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(wb_sel_i_3_bF_buf0_), .C(_37_), .Y(_38_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_38_), .C(_9__bF_buf6), .Y(_39_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_36_), .C(_39_), .Y(_2__30_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(ss_31_), .Y(_40_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf6_), .B(wb_dat_i[31]), .Y(_41_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(wb_sel_i_3_bF_buf5_), .C(_41_), .Y(_42_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_42_), .C(_9__bF_buf5), .Y(_43_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_40_), .C(_43_), .Y(_2__31_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(ss_16_), .Y(_44_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[16]), .B(wb_sel_i_2_bF_buf6_), .Y(_45_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(wb_sel_i_2_bF_buf5_), .C(_45_), .Y(_46_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_46_), .C(_9__bF_buf4), .Y(_47_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_44_), .C(_47_), .Y(_2__16_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(ss_17_), .Y(_48_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf4_), .B(wb_dat_i[17]), .Y(_49_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(wb_sel_i_2_bF_buf3_), .C(_49_), .Y(_50_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_50_), .C(_9__bF_buf3), .Y(_51_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_48_), .C(_51_), .Y(_2__17_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(ss_18_), .Y(_52_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf2_), .B(wb_dat_i[18]), .Y(_53_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(wb_sel_i_2_bF_buf1_), .C(_53_), .Y(_54_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_54_), .C(_9__bF_buf2), .Y(_55_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_52_), .C(_55_), .Y(_2__18_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(ss_19_), .Y(_56_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf0_), .B(wb_dat_i[19]), .Y(_57_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(wb_sel_i_2_bF_buf6_), .C(_57_), .Y(_58_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_58_), .C(_9__bF_buf1), .Y(_59_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_56_), .C(_59_), .Y(_2__19_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(ss_20_), .Y(_60_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf5_), .B(wb_dat_i[20]), .Y(_61_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(wb_sel_i_2_bF_buf4_), .C(_61_), .Y(_62_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_62_), .C(_9__bF_buf0), .Y(_63_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_60_), .C(_63_), .Y(_2__20_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(ss_21_), .Y(_64_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf3_), .B(wb_dat_i[21]), .Y(_65_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(wb_sel_i_2_bF_buf2_), .C(_65_), .Y(_66_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_66_), .C(_9__bF_buf6), .Y(_67_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_64_), .C(_67_), .Y(_2__21_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(ss_22_), .Y(_68_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf1_), .B(wb_dat_i[22]), .Y(_69_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(wb_sel_i_2_bF_buf0_), .C(_69_), .Y(_70_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_70_), .C(_9__bF_buf5), .Y(_71_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_68_), .C(_71_), .Y(_2__22_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(ss_23_), .Y(_72_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf6_), .B(wb_dat_i[23]), .Y(_73_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(wb_sel_i_2_bF_buf5_), .C(_73_), .Y(_74_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_74_), .C(_9__bF_buf4), .Y(_75_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_72_), .C(_75_), .Y(_2__23_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(ss_8_), .Y(_76_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[8]), .B(wb_sel_i_1_bF_buf7_), .Y(_77_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(wb_sel_i_1_bF_buf6_), .C(_77_), .Y(_78_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_78_), .C(_9__bF_buf3), .Y(_79_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_76_), .C(_79_), .Y(_2__8_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(ss_9_), .Y(_80_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf5_), .B(wb_dat_i[9]), .Y(_81_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(wb_sel_i_1_bF_buf4_), .C(_81_), .Y(_82_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_82_), .C(_9__bF_buf2), .Y(_83_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_80_), .C(_83_), .Y(_2__9_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(ss_10_), .Y(_84_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf3_), .B(wb_dat_i[10]), .Y(_85_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(wb_sel_i_1_bF_buf2_), .C(_85_), .Y(_86_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_86_), .C(_9__bF_buf1), .Y(_87_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_84_), .C(_87_), .Y(_2__10_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(ss_11_), .Y(_88_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf1_), .B(wb_dat_i[11]), .Y(_89_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(wb_sel_i_1_bF_buf0_), .C(_89_), .Y(_90_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_90_), .C(_9__bF_buf0), .Y(_91_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_88_), .C(_91_), .Y(_2__11_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(ss_12_), .Y(_92_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf7_), .B(wb_dat_i[12]), .Y(_93_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(wb_sel_i_1_bF_buf6_), .C(_93_), .Y(_94_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_94_), .C(_9__bF_buf6), .Y(_95_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_92_), .C(_95_), .Y(_2__12_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(ss_13_), .Y(_96_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf5_), .B(wb_dat_i[13]), .Y(_97_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(wb_sel_i_1_bF_buf4_), .C(_97_), .Y(_98_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_98_), .C(_9__bF_buf5), .Y(_99_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_96_), .C(_99_), .Y(_2__13_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(ss_14_), .Y(_100_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf3_), .B(wb_dat_i[14]), .Y(_101_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(wb_sel_i_1_bF_buf2_), .C(_101_), .Y(_102_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_102_), .C(_9__bF_buf4), .Y(_103_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_100_), .C(_103_), .Y(_2__14_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(ss_15_), .Y(_104_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf1_), .B(wb_dat_i[15]), .Y(_105_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(wb_sel_i_1_bF_buf0_), .C(_105_), .Y(_106_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_106_), .C(_9__bF_buf3), .Y(_107_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_104_), .C(_107_), .Y(_2__15_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(ss_0_), .Y(_108_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[0]), .B(wb_sel_i_0_bF_buf7_), .Y(_109_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(wb_sel_i_0_bF_buf6_), .C(_109_), .Y(_110_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_110_), .C(_9__bF_buf2), .Y(_111_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_108_), .C(_111_), .Y(_2__0_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(ss_1_), .Y(_112_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf5_), .B(wb_dat_i[1]), .Y(_113_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(wb_sel_i_0_bF_buf4_), .C(_113_), .Y(_114_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_114_), .C(_9__bF_buf1), .Y(_115_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_112_), .C(_115_), .Y(_2__1_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(ss_2_), .Y(_116_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf3_), .B(wb_dat_i[2]), .Y(_117_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(wb_sel_i_0_bF_buf2_), .C(_117_), .Y(_118_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_118_), .C(_9__bF_buf0), .Y(_119_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_116_), .C(_119_), .Y(_2__2_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(ss_3_), .Y(_120_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf1_), .B(wb_dat_i[3]), .Y(_121_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(wb_sel_i_0_bF_buf0_), .C(_121_), .Y(_122_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_122_), .C(_9__bF_buf6), .Y(_123_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf2), .B(_120_), .C(_123_), .Y(_2__3_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(ss_4_), .Y(_124_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf7_), .B(wb_dat_i[4]), .Y(_125_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(wb_sel_i_0_bF_buf6_), .C(_125_), .Y(_126_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_126_), .C(_9__bF_buf5), .Y(_127_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf1), .B(_124_), .C(_127_), .Y(_2__4_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(ss_5_), .Y(_128_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf5_), .B(wb_dat_i[5]), .Y(_129_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(wb_sel_i_0_bF_buf4_), .C(_129_), .Y(_130_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_130_), .C(_9__bF_buf4), .Y(_131_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf0), .B(_128_), .C(_131_), .Y(_2__5_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(ss_6_), .Y(_132_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf3_), .B(wb_dat_i[6]), .Y(_133_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(wb_sel_i_0_bF_buf2_), .C(_133_), .Y(_134_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_134_), .C(_9__bF_buf3), .Y(_135_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf4), .B(_132_), .C(_135_), .Y(_2__6_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(ss_7_), .Y(_136_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf1_), .B(wb_dat_i[7]), .Y(_137_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(wb_sel_i_0_bF_buf0_), .C(_137_), .Y(_138_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_138_), .C(_9__bF_buf2), .Y(_139_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_12__bF_buf3), .B(_136_), .C(_139_), .Y(_2__7_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .Y(_140_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[3]), .Y(_141_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[4]), .B(_7_), .C(_141_), .Y(_142_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_11__bF_buf6), .Y(_144_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(wb_sel_i_1_bF_buf7_), .C(_81_), .Y(_145_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_11__bF_buf5), .C(_143_), .Y(_146_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_140_), .C(_146_), .Y(_0__9_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(shift_tx_negedge), .Y(_147_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(wb_sel_i_1_bF_buf6_), .C(_85_), .Y(_148_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_11__bF_buf4), .C(_143_), .Y(_149_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_147_), .C(_149_), .Y(_0__10_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf3), .Y(_150_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(wb_sel_i_1_bF_buf5_), .C(_89_), .Y(_151_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_11__bF_buf3), .C(_143_), .Y(_152_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_150_), .C(_152_), .Y(_0__11_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(ie), .Y(_153_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(wb_sel_i_1_bF_buf4_), .C(_93_), .Y(_154_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_11__bF_buf2), .C(_143_), .Y(_155_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_153_), .C(_155_), .Y(_0__12_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(ass), .Y(_156_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(wb_sel_i_1_bF_buf3_), .C(_97_), .Y(_157_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_11__bF_buf1), .C(_143_), .Y(_158_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_156__bF_buf3), .C(_158_), .Y(_0__13_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(clgen_go), .Y(_159_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(wb_sel_i_1_bF_buf2_), .C(_77_), .Y(_160_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_11__bF_buf0), .C(_143_), .Y(_161_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf8), .B(clgen_last_clk), .C(clgen_pos_edge), .Y(_162_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(clgen_go), .B(_162_), .Y(_163_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_163_), .C(_161_), .Y(_0__8_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .Y(_164_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(wb_sel_i_0_bF_buf7_), .C(_109_), .Y(_165_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_11__bF_buf7), .C(_143_), .Y(_166_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_164_), .C(_166_), .Y(_0__0_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(char_len_1_), .Y(_167_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(wb_sel_i_0_bF_buf6_), .C(_113_), .Y(_168_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_11__bF_buf6), .C(_143_), .Y(_169_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_167_), .C(_169_), .Y(_0__1_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(char_len_2_), .Y(_170_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(wb_sel_i_0_bF_buf5_), .C(_117_), .Y(_171_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_11__bF_buf5), .C(_143_), .Y(_172_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_170_), .C(_172_), .Y(_0__2_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(char_len_3_), .Y(_173_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(wb_sel_i_0_bF_buf4_), .C(_121_), .Y(_174_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_11__bF_buf4), .C(_143_), .Y(_175_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_173_), .C(_175_), .Y(_0__3_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .Y(_176_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(wb_sel_i_0_bF_buf3_), .C(_125_), .Y(_177_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_11__bF_buf3), .C(_143_), .Y(_178_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_176_), .C(_178_), .Y(_0__4_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .Y(_179_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(wb_sel_i_0_bF_buf2_), .C(_129_), .Y(_180_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_11__bF_buf2), .C(_143_), .Y(_181_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_179_), .C(_181_), .Y(_0__5_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(char_len_6_), .Y(_182_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(wb_sel_i_0_bF_buf1_), .C(_133_), .Y(_183_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_11__bF_buf1), .C(_143_), .Y(_184_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_182_), .C(_184_), .Y(_0__6_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(ctrl_7_), .Y(_185_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(wb_sel_i_0_bF_buf0_), .C(_137_), .Y(_186_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_11__bF_buf0), .C(_143_), .Y(_187_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_185_), .C(_187_), .Y(_0__7_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_8_), .Y(_188_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[4]), .B(wb_adr_i[2]), .C(_141_), .Y(_189_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(_189__bF_buf3), .Y(_190_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_190__bF_buf3), .B(_11__bF_buf7), .Y(_191_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(wb_sel_i_1_bF_buf1_), .C(_77_), .Y(_192_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_192_), .C(_190__bF_buf2), .Y(_193_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_188_), .C(_193_), .Y(_1__8_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_9_), .Y(_194_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(wb_sel_i_1_bF_buf0_), .C(_81_), .Y(_195_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_195_), .C(_190__bF_buf1), .Y(_196_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_194_), .C(_196_), .Y(_1__9_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_10_), .Y(_197_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(wb_sel_i_1_bF_buf7_), .C(_85_), .Y(_198_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_198_), .C(_190__bF_buf0), .Y(_199_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_197_), .C(_199_), .Y(_1__10_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_11_), .Y(_200_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(wb_sel_i_1_bF_buf6_), .C(_89_), .Y(_201_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_201_), .C(_190__bF_buf3), .Y(_202_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_200_), .C(_202_), .Y(_1__11_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_12_), .Y(_203_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(wb_sel_i_1_bF_buf5_), .C(_93_), .Y(_204_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_204_), .C(_190__bF_buf2), .Y(_205_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_203_), .C(_205_), .Y(_1__12_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_13_), .Y(_206_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(wb_sel_i_1_bF_buf4_), .C(_97_), .Y(_207_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_207_), .C(_190__bF_buf1), .Y(_208_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_206_), .C(_208_), .Y(_1__13_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_14_), .Y(_209_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(wb_sel_i_1_bF_buf3_), .C(_101_), .Y(_210_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_210_), .C(_190__bF_buf0), .Y(_211_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_209_), .C(_211_), .Y(_1__14_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_15_), .Y(_212_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(wb_sel_i_1_bF_buf2_), .C(_105_), .Y(_213_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_213_), .C(_190__bF_buf3), .Y(_214_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_212_), .C(_214_), .Y(_1__15_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_0_), .Y(_215_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(wb_sel_i_0_bF_buf7_), .C(_109_), .Y(_216_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf6), .B(_216_), .C(_190__bF_buf2), .Y(_217_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_215_), .C(_217_), .Y(_1__0_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_1_), .Y(_218_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(wb_sel_i_0_bF_buf6_), .C(_113_), .Y(_219_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf5), .B(_219_), .C(_190__bF_buf1), .Y(_220_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_218_), .C(_220_), .Y(_1__1_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_2_), .Y(_221_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(wb_sel_i_0_bF_buf5_), .C(_117_), .Y(_222_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf4), .B(_222_), .C(_190__bF_buf0), .Y(_223_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_221_), .C(_223_), .Y(_1__2_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_3_), .Y(_224_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(wb_sel_i_0_bF_buf4_), .C(_121_), .Y(_225_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf3), .B(_225_), .C(_190__bF_buf3), .Y(_226_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_224_), .C(_226_), .Y(_1__3_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_4_), .Y(_227_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(wb_sel_i_0_bF_buf3_), .C(_125_), .Y(_228_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf2), .B(_228_), .C(_190__bF_buf2), .Y(_229_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_227_), .C(_229_), .Y(_1__4_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_5_), .Y(_230_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(wb_sel_i_0_bF_buf2_), .C(_129_), .Y(_231_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf1), .B(_231_), .C(_190__bF_buf1), .Y(_232_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_230_), .C(_232_), .Y(_1__5_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_6_), .Y(_233_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(wb_sel_i_0_bF_buf1_), .C(_133_), .Y(_234_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf0), .B(_234_), .C(_190__bF_buf0), .Y(_235_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_233_), .C(_235_), .Y(_1__6_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_7_), .Y(_236_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(wb_sel_i_0_bF_buf0_), .C(_137_), .Y(_237_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_11__bF_buf7), .B(_237_), .C(_190__bF_buf3), .Y(_238_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_236_), .C(_238_), .Y(_1__7_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(rx_64_), .Y(_239_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(rx_32_), .Y(_240_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[4]), .Y(_241_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[2]), .B(_241_), .C(_141_), .Y(_242_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[3]), .B(_241_), .C(_7_), .Y(_243_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf3), .B(_240_), .C(_239_), .D(_243__bF_buf3), .Y(_244_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf2), .B(_108_), .C(_215_), .D(_189__bF_buf2), .Y(_245_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_244_), .Y(_246_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_7_), .C(_141_), .Y(_247_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[2]), .B(wb_adr_i[3]), .Y(_248_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_248_), .C(_247_), .Y(_249_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(rx_96_), .Y(_250_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(wb_adr_i[2]), .B(wb_adr_i[3]), .C(_241_), .Y(_251_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_250_), .C(_142_), .D(_164_), .Y(_252_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_0_), .B(_249__bF_buf4), .C(_252_), .Y(_253_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_246_), .Y(wb_dat_0_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(rx_65_), .Y(_254_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(rx_33_), .Y(_255_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf2), .B(_255_), .C(_254_), .D(_243__bF_buf2), .Y(_256_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf1), .B(_112_), .C(_218_), .D(_189__bF_buf1), .Y(_257_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_256_), .Y(_258_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(rx_97_), .Y(_259_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_259_), .C(_142_), .D(_167_), .Y(_260_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(rx_1_), .B(_249__bF_buf3), .C(_260_), .Y(_261_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_258_), .Y(wb_dat_1_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(rx_66_), .Y(_262_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(rx_34_), .Y(_263_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf1), .B(_263_), .C(_262_), .D(_243__bF_buf1), .Y(_264_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf0), .B(_116_), .C(_221_), .D(_189__bF_buf0), .Y(_265_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_264_), .Y(_266_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(rx_98_), .Y(_267_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_267_), .C(_142_), .D(_170_), .Y(_268_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(rx_2_), .B(_249__bF_buf2), .C(_268_), .Y(_269_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_266_), .Y(wb_dat_2_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(rx_67_), .Y(_270_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(rx_35_), .Y(_271_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf0), .B(_271_), .C(_270_), .D(_243__bF_buf0), .Y(_272_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf3), .B(_120_), .C(_224_), .D(_189__bF_buf3), .Y(_273_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_272_), .Y(_274_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(rx_99_), .Y(_275_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_275_), .C(_142_), .D(_173_), .Y(_276_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(rx_3_), .B(_249__bF_buf1), .C(_276_), .Y(_277_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_274_), .Y(wb_dat_3_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(rx_68_), .Y(_278_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(rx_36_), .Y(_279_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf3), .B(_279_), .C(_278_), .D(_243__bF_buf3), .Y(_280_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf2), .B(_124_), .C(_227_), .D(_189__bF_buf2), .Y(_281_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_280_), .Y(_282_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(rx_100_), .Y(_283_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_283_), .C(_142_), .D(_176_), .Y(_284_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(rx_4_), .B(_249__bF_buf0), .C(_284_), .Y(_285_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_282_), .Y(wb_dat_4_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf1), .B(_128_), .C(_230_), .D(_189__bF_buf1), .Y(_286_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(rx_69_), .Y(_287_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(rx_37_), .Y(_288_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf2), .B(_288_), .C(_287_), .D(_243__bF_buf2), .Y(_289_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_289_), .Y(_290_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(rx_101_), .Y(_291_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_291_), .C(_142_), .D(_179_), .Y(_292_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(rx_5_), .B(_249__bF_buf4), .C(_292_), .Y(_293_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_290_), .Y(wb_dat_5_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(rx_70_), .Y(_294_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(rx_38_), .Y(_295_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf1), .B(_295_), .C(_294_), .D(_243__bF_buf1), .Y(_296_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf0), .B(_132_), .C(_233_), .D(_189__bF_buf0), .Y(_297_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_296_), .Y(_298_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(rx_102_), .Y(_299_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_299_), .C(_142_), .D(_182_), .Y(_300_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(rx_6_), .B(_249__bF_buf3), .C(_300_), .Y(_301_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_298_), .Y(wb_dat_6_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(rx_71_), .Y(_302_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(rx_39_), .Y(_303_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf0), .B(_303_), .C(_302_), .D(_243__bF_buf0), .Y(_304_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf3), .B(_136_), .C(_236_), .D(_189__bF_buf3), .Y(_305_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_304_), .Y(_306_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(rx_103_), .Y(_307_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_307_), .C(_142_), .D(_185_), .Y(_308_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(rx_7_), .B(_249__bF_buf2), .C(_308_), .Y(_309_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_306_), .Y(wb_dat_7_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(rx_72_), .Y(_310_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(rx_40_), .Y(_311_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf3), .B(_311_), .C(_310_), .D(_243__bF_buf3), .Y(_312_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf2), .B(_76_), .C(_188_), .D(_189__bF_buf2), .Y(_313_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_312_), .Y(_314_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(rx_104_), .Y(_315_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_315_), .C(_142_), .D(_159_), .Y(_316_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(rx_8_), .B(_249__bF_buf1), .C(_316_), .Y(_317_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_314_), .Y(wb_dat_8_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(rx_73_), .Y(_318_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(rx_41_), .Y(_319_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf2), .B(_319_), .C(_318_), .D(_243__bF_buf2), .Y(_320_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf1), .B(_80_), .C(_194_), .D(_189__bF_buf1), .Y(_321_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_320_), .Y(_322_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(rx_105_), .Y(_323_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_323_), .C(_142_), .D(_140_), .Y(_324_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(rx_9_), .B(_249__bF_buf0), .C(_324_), .Y(_325_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_322_), .Y(wb_dat_9_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(rx_74_), .Y(_326_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(rx_42_), .Y(_327_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf1), .B(_327_), .C(_326_), .D(_243__bF_buf1), .Y(_328_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf0), .B(_84_), .C(_197_), .D(_189__bF_buf0), .Y(_329_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_328_), .Y(_330_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(rx_106_), .Y(_331_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_331_), .C(_142_), .D(_147_), .Y(_332_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(rx_10_), .B(_249__bF_buf4), .C(_332_), .Y(_333_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_330_), .Y(wb_dat_10_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(rx_75_), .Y(_334_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(rx_43_), .Y(_335_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf0), .B(_335_), .C(_334_), .D(_243__bF_buf0), .Y(_336_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf3), .B(_88_), .C(_200_), .D(_189__bF_buf3), .Y(_337_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_336_), .Y(_338_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(rx_107_), .Y(_339_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_339_), .C(_142_), .D(_150_), .Y(_340_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(rx_11_), .B(_249__bF_buf3), .C(_340_), .Y(_341_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_338_), .Y(wb_dat_11_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(rx_76_), .Y(_342_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(rx_44_), .Y(_343_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf3), .B(_343_), .C(_342_), .D(_243__bF_buf3), .Y(_344_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf2), .B(_92_), .C(_203_), .D(_189__bF_buf2), .Y(_345_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_344_), .Y(_346_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(rx_108_), .Y(_347_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_347_), .C(_142_), .D(_153_), .Y(_348_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(rx_12_), .B(_249__bF_buf2), .C(_348_), .Y(_349_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_346_), .Y(wb_dat_12_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf1), .B(_96_), .C(_206_), .D(_189__bF_buf1), .Y(_350_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(rx_77_), .Y(_351_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(rx_45_), .Y(_352_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf2), .B(_352_), .C(_351_), .D(_243__bF_buf2), .Y(_353_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_353_), .Y(_354_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(rx_109_), .Y(_355_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_355_), .C(_142_), .D(_156__bF_buf2), .Y(_356_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(rx_13_), .B(_249__bF_buf1), .C(_356_), .Y(_357_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_354_), .Y(wb_dat_13_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(_251_), .Y(_358_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(rx_46_), .Y(_359_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_189__bF_buf0), .B(_209_), .C(_242__bF_buf1), .D(_359_), .Y(_360_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(rx_110_), .B(_358__bF_buf3), .C(_360_), .Y(_361_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(rx_78_), .Y(_362_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf0), .B(_100_), .C(_243__bF_buf1), .D(_362_), .Y(_363_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(rx_14_), .B(_249__bF_buf0), .C(_363_), .Y(_364_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_364_), .Y(wb_dat_14_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(rx_47_), .Y(_365_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_189__bF_buf3), .B(_212_), .C(_242__bF_buf0), .D(_365_), .Y(_366_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(rx_111_), .B(_358__bF_buf2), .C(_366_), .Y(_367_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(rx_79_), .Y(_368_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_8__bF_buf3), .B(_104_), .C(_243__bF_buf0), .D(_368_), .Y(_369_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(rx_15_), .B(_249__bF_buf4), .C(_369_), .Y(_370_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_370_), .Y(wb_dat_15_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(rx_16_), .B(_249__bF_buf3), .Y(_371_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(_242__bF_buf3), .Y(_372_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(_243__bF_buf3), .Y(_373_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_48_), .C(rx_80_), .D(_373_), .Y(_374_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf1), .B(ss_16_), .C(rx_112_), .D(_358__bF_buf1), .Y(_375_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_375_), .C(_374_), .Y(wb_dat_16_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(rx_17_), .B(_249__bF_buf2), .Y(_376_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_49_), .C(rx_81_), .D(_373_), .Y(_377_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf0), .B(ss_17_), .C(rx_113_), .D(_358__bF_buf0), .Y(_378_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_378_), .C(_377_), .Y(wb_dat_17_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(rx_18_), .B(_249__bF_buf1), .Y(_379_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_50_), .C(rx_82_), .D(_373_), .Y(_380_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf6), .B(ss_18_), .C(rx_114_), .D(_358__bF_buf3), .Y(_381_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_381_), .C(_380_), .Y(wb_dat_18_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(rx_19_), .B(_249__bF_buf0), .Y(_382_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_51_), .C(rx_83_), .D(_373_), .Y(_383_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf5), .B(ss_19_), .C(rx_115_), .D(_358__bF_buf2), .Y(_384_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_384_), .C(_383_), .Y(wb_dat_19_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(rx_20_), .B(_249__bF_buf4), .Y(_385_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_52_), .C(rx_84_), .D(_373_), .Y(_386_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf4), .B(ss_20_), .C(rx_116_), .D(_358__bF_buf1), .Y(_387_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_387_), .C(_386_), .Y(wb_dat_20_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(rx_21_), .B(_249__bF_buf3), .Y(_388_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_53_), .C(rx_85_), .D(_373_), .Y(_389_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf3), .B(ss_21_), .C(rx_117_), .D(_358__bF_buf0), .Y(_390_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_390_), .C(_389_), .Y(wb_dat_21_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(rx_22_), .B(_249__bF_buf2), .Y(_391_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_54_), .C(rx_86_), .D(_373_), .Y(_392_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf2), .B(ss_22_), .C(rx_118_), .D(_358__bF_buf3), .Y(_393_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(wb_dat_22_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(rx_23_), .B(_249__bF_buf1), .Y(_394_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_55_), .C(rx_87_), .D(_373_), .Y(_395_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf1), .B(ss_23_), .C(rx_119_), .D(_358__bF_buf2), .Y(_396_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_396_), .C(_395_), .Y(wb_dat_23_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(rx_24_), .B(_249__bF_buf0), .Y(_397_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_56_), .C(rx_88_), .D(_373_), .Y(_398_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf0), .B(ss_24_), .C(rx_120_), .D(_358__bF_buf1), .Y(_399_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_399_), .C(_398_), .Y(wb_dat_24_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(rx_25_), .B(_249__bF_buf4), .Y(_400_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_57_), .C(rx_89_), .D(_373_), .Y(_401_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf6), .B(ss_25_), .C(rx_121_), .D(_358__bF_buf0), .Y(_402_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_402_), .C(_401_), .Y(wb_dat_25_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(rx_26_), .B(_249__bF_buf3), .Y(_403_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_58_), .C(rx_90_), .D(_373_), .Y(_404_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf5), .B(ss_26_), .C(rx_122_), .D(_358__bF_buf3), .Y(_405_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_404_), .Y(wb_dat_26_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(rx_27_), .B(_249__bF_buf2), .Y(_406_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_59_), .C(rx_91_), .D(_373_), .Y(_407_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf4), .B(ss_27_), .C(rx_123_), .D(_358__bF_buf2), .Y(_408_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_408_), .C(_407_), .Y(wb_dat_27_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(rx_28_), .B(_249__bF_buf1), .Y(_409_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_60_), .C(rx_92_), .D(_373_), .Y(_410_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf3), .B(ss_28_), .C(rx_124_), .D(_358__bF_buf1), .Y(_411_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_411_), .C(_410_), .Y(wb_dat_28_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(rx_29_), .B(_249__bF_buf0), .Y(_412_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_61_), .C(rx_93_), .D(_373_), .Y(_413_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf2), .B(ss_29_), .C(rx_125_), .D(_358__bF_buf0), .Y(_414_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(wb_dat_29_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(rx_30_), .B(_249__bF_buf4), .Y(_415_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_62_), .C(rx_94_), .D(_373_), .Y(_416_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf1), .B(ss_30_), .C(rx_126_), .D(_358__bF_buf3), .Y(_417_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_417_), .C(_416_), .Y(wb_dat_30_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(rx_31_), .B(_249__bF_buf3), .Y(_418_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(rx_63_), .C(rx_95_), .D(_373_), .Y(_419_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_9__bF_buf0), .B(ss_31_), .C(rx_127_), .D(_358__bF_buf2), .Y(_420_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_420_), .C(_419_), .Y(wb_dat_31_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf7), .C(ss_0_), .Y(_425__0_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf6), .C(ss_1_), .Y(_425__1_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf5), .C(ss_2_), .Y(_425__2_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf4), .C(ss_3_), .Y(_425__3_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf3), .C(ss_4_), .Y(_425__4_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf2), .C(ss_5_), .Y(_425__5_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf1), .C(ss_6_), .Y(_425__6_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf0), .C(ss_7_), .Y(_425__7_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf9), .C(ss_8_), .Y(_425__8_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf8), .C(ss_9_), .Y(_425__9_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf7), .C(ss_10_), .Y(_425__10_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf6), .C(ss_11_), .Y(_425__11_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf5), .C(ss_12_), .Y(_425__12_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf4), .C(ss_13_), .Y(_425__13_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf3), .C(ss_14_), .Y(_425__14_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf2), .C(ss_15_), .Y(_425__15_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf1), .C(ss_16_), .Y(_425__16_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf0), .C(ss_17_), .Y(_425__17_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf9), .C(ss_18_), .Y(_425__18_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf8), .C(ss_19_), .Y(_425__19_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf7), .C(ss_20_), .Y(_425__20_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf6), .C(ss_21_), .Y(_425__21_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf5), .C(ss_22_), .Y(_425__22_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf4), .C(ss_23_), .Y(_425__23_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf3), .C(ss_24_), .Y(_425__24_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf2), .C(ss_25_), .Y(_425__25_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf1), .C(ss_26_), .Y(_425__26_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(clgen_enable_bF_buf0), .C(ss_27_), .Y(_425__27_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(clgen_enable_bF_buf9), .C(ss_28_), .Y(_425__28_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(clgen_enable_bF_buf8), .C(ss_29_), .Y(_425__29_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf1), .B(clgen_enable_bF_buf7), .C(ss_30_), .Y(_425__30_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(clgen_enable_bF_buf6), .C(ss_31_), .Y(_425__31_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(wb_stb_i), .B(wb_cyc_i), .Y(_421_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_421_), .Y(_3_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_247_), .Y(shift_latch_0_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_242__bF_buf2), .Y(shift_latch_1_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_243__bF_buf2), .Y(shift_latch_2_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_251_), .Y(shift_latch_3_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(_422_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_422_), .C(_162_), .D(_153_), .Y(_4_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(wb_rst_i), .Y(_5_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_423_), .Y(mosi_pad_o) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_424_), .Y(sclk_pad_o) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_425__0_), .Y(ss_pad_o[0]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_425__1_), .Y(ss_pad_o[1]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_425__2_), .Y(ss_pad_o[2]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_425__3_), .Y(ss_pad_o[3]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_425__4_), .Y(ss_pad_o[4]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_425__5_), .Y(ss_pad_o[5]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_425__6_), .Y(ss_pad_o[6]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_425__7_), .Y(ss_pad_o[7]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_425__8_), .Y(ss_pad_o[8]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_425__9_), .Y(ss_pad_o[9]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_425__10_), .Y(ss_pad_o[10]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_425__11_), .Y(ss_pad_o[11]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_425__12_), .Y(ss_pad_o[12]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_425__13_), .Y(ss_pad_o[13]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_425__14_), .Y(ss_pad_o[14]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_425__15_), .Y(ss_pad_o[15]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_425__16_), .Y(ss_pad_o[16]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_425__17_), .Y(ss_pad_o[17]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_425__18_), .Y(ss_pad_o[18]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_425__19_), .Y(ss_pad_o[19]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_425__20_), .Y(ss_pad_o[20]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_425__21_), .Y(ss_pad_o[21]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_425__22_), .Y(ss_pad_o[22]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_425__23_), .Y(ss_pad_o[23]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_425__24_), .Y(ss_pad_o[24]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_425__25_), .Y(ss_pad_o[25]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_425__26_), .Y(ss_pad_o[26]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_425__27_), .Y(ss_pad_o[27]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_425__28_), .Y(ss_pad_o[28]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_425__29_), .Y(ss_pad_o[29]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_425__30_), .Y(ss_pad_o[30]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_425__31_), .Y(ss_pad_o[31]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_426_), .Y(wb_ack_o) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_427__0_), .Y(wb_dat_o[0]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_427__1_), .Y(wb_dat_o[1]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_427__2_), .Y(wb_dat_o[2]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_427__3_), .Y(wb_dat_o[3]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_427__4_), .Y(wb_dat_o[4]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_427__5_), .Y(wb_dat_o[5]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_427__6_), .Y(wb_dat_o[6]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_427__7_), .Y(wb_dat_o[7]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_427__8_), .Y(wb_dat_o[8]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_427__9_), .Y(wb_dat_o[9]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_427__10_), .Y(wb_dat_o[10]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_427__11_), .Y(wb_dat_o[11]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_427__12_), .Y(wb_dat_o[12]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_427__13_), .Y(wb_dat_o[13]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_427__14_), .Y(wb_dat_o[14]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_427__15_), .Y(wb_dat_o[15]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_427__16_), .Y(wb_dat_o[16]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_427__17_), .Y(wb_dat_o[17]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_427__18_), .Y(wb_dat_o[18]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_427__19_), .Y(wb_dat_o[19]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_427__20_), .Y(wb_dat_o[20]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_427__21_), .Y(wb_dat_o[21]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_427__22_), .Y(wb_dat_o[22]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_427__23_), .Y(wb_dat_o[23]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_427__24_), .Y(wb_dat_o[24]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_427__25_), .Y(wb_dat_o[25]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_427__26_), .Y(wb_dat_o[26]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_427__27_), .Y(wb_dat_o[27]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_427__28_), .Y(wb_dat_o[28]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_427__29_), .Y(wb_dat_o[29]) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_427__30_), .Y(wb_dat_o[30]) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_427__31_), .Y(wb_dat_o[31]) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(wb_err_o) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(wb_int_o) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf3), .D(_2__0_), .Q(ss_0_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf3), .D(_2__1_), .Q(ss_1_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf3), .D(_2__2_), .Q(ss_2_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf3), .D(_2__3_), .Q(ss_3_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf3), .D(_2__4_), .Q(ss_4_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf3), .D(_2__5_), .Q(ss_5_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf3), .D(_2__6_), .Q(ss_6_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf3), .D(_2__7_), .Q(ss_7_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf3), .D(_2__8_), .Q(ss_8_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf3), .D(_2__9_), .Q(ss_9_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf3), .D(_2__10_), .Q(ss_10_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf3), .D(_2__11_), .Q(ss_11_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf3), .D(_2__12_), .Q(ss_12_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_2__13_), .Q(ss_13_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_2__14_), .Q(ss_14_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf2), .D(_2__15_), .Q(ss_15_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf2), .D(_2__16_), .Q(ss_16_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf2), .D(_2__17_), .Q(ss_17_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf2), .D(_2__18_), .Q(ss_18_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf2), .D(_2__19_), .Q(ss_19_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf2), .D(_2__20_), .Q(ss_20_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf2), .D(_2__21_), .Q(ss_21_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf2), .D(_2__22_), .Q(ss_22_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf2), .D(_2__23_), .Q(ss_23_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf2), .D(_2__24_), .Q(ss_24_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf2), .D(_2__25_), .Q(ss_25_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf2), .D(_2__26_), .Q(ss_26_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf2), .D(_2__27_), .Q(ss_27_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_2__28_), .Q(ss_28_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_2__29_), .Q(ss_29_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf1), .D(_2__30_), .Q(ss_30_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf1), .D(_2__31_), .Q(ss_31_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf1), .D(_0__0_), .Q(char_len_0_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf1), .D(_0__1_), .Q(char_len_1_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf1), .D(_0__2_), .Q(char_len_2_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf1), .D(_0__3_), .Q(char_len_3_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf1), .D(_0__4_), .Q(char_len_4_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_38 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf1), .D(_0__5_), .Q(char_len_5_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_39 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf1), .D(_0__6_), .Q(char_len_6_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_40 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf1), .D(_0__7_), .Q(ctrl_7_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_41 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf1), .D(_0__8_), .Q(clgen_go), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_42 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf1), .D(_0__9_), .Q(rx_negedge), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_43 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf1), .D(_0__10_), .Q(shift_tx_negedge), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_44 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_0__11_), .Q(lsb), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_45 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_0__12_), .Q(ie), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_46 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf0), .D(_0__13_), .Q(ass), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_47 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf0), .D(_1__0_), .Q(clgen_divider_0_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_48 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf0), .D(_1__1_), .Q(clgen_divider_1_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_49 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf0), .D(_1__2_), .Q(clgen_divider_2_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_50 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf0), .D(_1__3_), .Q(clgen_divider_3_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_51 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf0), .D(_1__4_), .Q(clgen_divider_4_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_52 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf0), .D(_1__5_), .Q(clgen_divider_5_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_53 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf0), .D(_1__6_), .Q(clgen_divider_6_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_54 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf0), .D(_1__7_), .Q(clgen_divider_7_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_55 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf0), .D(_1__8_), .Q(clgen_divider_8_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_56 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf0), .D(_1__9_), .Q(clgen_divider_9_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_57 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf0), .D(_1__10_), .Q(clgen_divider_10_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_58 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf0), .D(_1__11_), .Q(clgen_divider_11_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_59 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_1__12_), .Q(clgen_divider_12_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_60 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_1__13_), .Q(clgen_divider_13_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_61 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf3), .D(_1__14_), .Q(clgen_divider_14_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_62 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf3), .D(_1__15_), .Q(clgen_divider_15_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_63 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf3), .D(_4_), .Q(_428_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_64 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf3), .D(_3_), .Q(_426_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_65 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf3), .D(wb_dat_0_), .Q(_427__0_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_66 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf3), .D(wb_dat_1_), .Q(_427__1_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_67 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf3), .D(wb_dat_2_), .Q(_427__2_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_68 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf3), .D(wb_dat_3_), .Q(_427__3_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_69 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf3), .D(wb_dat_4_), .Q(_427__4_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_70 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf3), .D(wb_dat_5_), .Q(_427__5_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_71 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf3), .D(wb_dat_6_), .Q(_427__6_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_72 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf3), .D(wb_dat_7_), .Q(_427__7_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_73 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf3), .D(wb_dat_8_), .Q(_427__8_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_74 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(wb_dat_9_), .Q(_427__9_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_75 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(wb_dat_10_), .Q(_427__10_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_76 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf2), .D(wb_dat_11_), .Q(_427__11_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_77 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf2), .D(wb_dat_12_), .Q(_427__12_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_78 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf2), .D(wb_dat_13_), .Q(_427__13_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_79 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf2), .D(wb_dat_14_), .Q(_427__14_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_80 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf2), .D(wb_dat_15_), .Q(_427__15_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_81 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf2), .D(wb_dat_16_), .Q(_427__16_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_82 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf2), .D(wb_dat_17_), .Q(_427__17_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_83 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf2), .D(wb_dat_18_), .Q(_427__18_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_84 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf2), .D(wb_dat_19_), .Q(_427__19_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_85 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf2), .D(wb_dat_20_), .Q(_427__20_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_86 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf2), .D(wb_dat_21_), .Q(_427__21_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_87 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf2), .D(wb_dat_22_), .Q(_427__22_), .R(_5__bF_buf3), .S(vdd) );
DFFSR DFFSR_88 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf2), .D(wb_dat_23_), .Q(_427__23_), .R(_5__bF_buf2), .S(vdd) );
DFFSR DFFSR_89 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(wb_dat_24_), .Q(_427__24_), .R(_5__bF_buf1), .S(vdd) );
DFFSR DFFSR_90 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(wb_dat_25_), .Q(_427__25_), .R(_5__bF_buf0), .S(vdd) );
DFFSR DFFSR_91 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf1), .D(wb_dat_26_), .Q(_427__26_), .R(_5__bF_buf8), .S(vdd) );
DFFSR DFFSR_92 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf1), .D(wb_dat_27_), .Q(_427__27_), .R(_5__bF_buf7), .S(vdd) );
DFFSR DFFSR_93 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf1), .D(wb_dat_28_), .Q(_427__28_), .R(_5__bF_buf6), .S(vdd) );
DFFSR DFFSR_94 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf1), .D(wb_dat_29_), .Q(_427__29_), .R(_5__bF_buf5), .S(vdd) );
DFFSR DFFSR_95 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf1), .D(wb_dat_30_), .Q(_427__30_), .R(_5__bF_buf4), .S(vdd) );
DFFSR DFFSR_96 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf1), .D(wb_dat_31_), .Q(_427__31_), .R(_5__bF_buf3), .S(vdd) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf5), .Y(_503_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_424_), .Y(_504_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_9_), .B(clgen_cnt_10_), .Y(_505_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_11_), .B(clgen_cnt_12_), .Y(_506_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_506_), .Y(_507_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_13_), .B(clgen_cnt_14_), .Y(_508_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_8_), .B(clgen_cnt_15_), .Y(_509_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_509_), .Y(_510_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_510_), .Y(_511_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_4_), .B(clgen_cnt_7_), .Y(_512_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_5_), .B(clgen_cnt_6_), .Y(_513_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .Y(_514_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_1_), .Y(_515_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_3_), .B(clgen_cnt_2_), .Y(_516_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_0_), .B(_515_), .C(_516_), .Y(_517_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_517_), .Y(_518_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_518_), .Y(_519_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_15_), .Y(_520_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_12_), .Y(_521_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_521_), .Y(_522_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_10_), .B(clgen_divider_11_), .Y(_523_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_8_), .B(clgen_divider_9_), .Y(_524_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_14_), .B(clgen_divider_13_), .Y(_525_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_524_), .C(_525_), .Y(_526_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_526_), .Y(_527_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_2_), .B(clgen_divider_3_), .Y(_528_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_0_), .B(clgen_divider_1_), .Y(_529_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_529_), .Y(_530_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_6_), .B(clgen_divider_7_), .Y(_531_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_4_), .B(clgen_divider_5_), .Y(_532_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_532_), .Y(_533_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_533_), .Y(_534_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_527_), .Y(_535_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(clgen_go), .B(_503_), .C(_424_), .Y(_536_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_519_), .C(_535_), .D(_536_), .Y(_432_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf4), .B(_424_), .Y(_537_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_537_), .C(_535_), .D(_504_), .Y(_431_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_510_), .Y(_538_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .Y(_539_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_0_), .B(clgen_cnt_1_), .Y(_540_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_540_), .Y(_541_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_541_), .Y(_542_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_542_), .C(clgen_enable_bF_buf3), .Y(_434_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_540_), .Y(_435_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_435_), .Y(_436_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_511_), .Y(_437_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_437_), .Y(_438_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_0_), .Y(_439_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_0_), .B(_434_), .C(_439_), .Y(_430__0_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_0_), .B(clgen_cnt_1_), .Y(_440_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_1_), .Y(_441_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_440_), .C(_441_), .Y(_430__1_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_2_), .Y(_442_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_540_), .Y(_443_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_0_), .B(clgen_cnt_1_), .C(clgen_cnt_2_), .Y(_444_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_444_), .Y(_445_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_2_), .Y(_446_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_445_), .C(_446_), .Y(_430__2_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_3_), .B(_443_), .C(_541_), .Y(_447_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_3_), .Y(_448_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_447_), .C(_448_), .Y(_430__3_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_4_), .Y(_449_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_511_), .C(_503_), .Y(_450_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_4_), .B(_435_), .Y(_451_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_4_), .Y(_452_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_541_), .Y(_453_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_453_), .C(_450_), .Y(_454_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(_454_), .Y(_430__4_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(clgen_cnt_5_), .Y(_455_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_5_), .Y(_456_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_455_), .C(_456_), .Y(_430__5_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_451_), .Y(_457_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_541_), .Y(_458_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(clgen_cnt_5_), .C(clgen_cnt_6_), .Y(_459_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_457_), .Y(_460_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_6_), .Y(_461_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_434_), .C(_461_), .Y(_430__6_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_7_), .B(_457_), .C(_436_), .Y(_462_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_7_), .Y(_463_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_462_), .C(_463_), .Y(_430__7_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_8_), .Y(_464_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_8_), .Y(_465_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_436_), .Y(_466_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(clgen_cnt_8_), .C(_435_), .Y(_467_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_467_), .C(_450_), .Y(_468_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_450_), .C(_468_), .Y(_430__8_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_9_), .Y(_469_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_539_), .C(_541_), .Y(_470_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_469_), .Y(_471_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_9_), .Y(_472_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_434_), .C(_472_), .Y(_430__9_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_10_), .Y(_473_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_10_), .Y(_474_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_467_), .C(_474_), .Y(_475_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_505_), .Y(_476_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_470_), .Y(_477_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_450_), .Y(_478_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_450_), .C(_478_), .Y(_430__10_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_11_), .Y(_479_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_467_), .C(_479_), .Y(_480_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_11_), .B(_476_), .C(_470_), .Y(_481_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_480_), .C(_450_), .Y(_482_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_11_), .Y(_483_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_482_), .Y(_430__11_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_467_), .Y(_484_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(clgen_cnt_11_), .C(clgen_cnt_12_), .Y(_485_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_470_), .Y(_486_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_434_), .Y(_487_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_434_), .C(_487_), .D(_485_), .Y(_430__12_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_13_), .Y(_488_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_507_), .Y(_489_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_467_), .C(_488_), .Y(_490_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_13_), .B(_507_), .C(_470_), .Y(_491_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_490_), .C(_450_), .Y(_492_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_503_), .C(clgen_divider_13_), .Y(_493_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_492_), .Y(_430__13_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_467_), .Y(_494_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(clgen_cnt_13_), .C(clgen_cnt_14_), .Y(_495_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_486_), .C(_434_), .Y(_496_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(clgen_divider_14_), .B(_450_), .Y(_497_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_496_), .C(_497_), .Y(_430__14_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(clgen_cnt_15_), .Y(_498_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_508_), .Y(_499_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_499_), .C(_450_), .Y(_500_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_450_), .C(_500_), .D(_498_), .Y(_430__15_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_503_), .C(_424_), .Y(_501_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(clgen_last_clk), .Y(_502_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_502_), .C(_501_), .Y(_429_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(wb_rst_i), .Y(_433_) );
DFFSR DFFSR_97 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf1), .D(_432_), .Q(clgen_pos_edge), .R(_433__bF_buf3), .S(vdd) );
DFFSR DFFSR_98 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf1), .D(_431_), .Q(clgen_neg_edge), .R(_433__bF_buf2), .S(vdd) );
DFFSR DFFSR_99 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf1), .D(_429_), .Q(_424_), .R(_433__bF_buf1), .S(vdd) );
DFFSR DFFSR_100 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf1), .D(_430__0_), .Q(clgen_cnt_0_), .R(vdd), .S(_433__bF_buf0) );
DFFSR DFFSR_101 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf1), .D(_430__1_), .Q(clgen_cnt_1_), .R(vdd), .S(_433__bF_buf3) );
DFFSR DFFSR_102 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf1), .D(_430__2_), .Q(clgen_cnt_2_), .R(vdd), .S(_433__bF_buf2) );
DFFSR DFFSR_103 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf1), .D(_430__3_), .Q(clgen_cnt_3_), .R(vdd), .S(_433__bF_buf1) );
DFFSR DFFSR_104 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_430__4_), .Q(clgen_cnt_4_), .R(vdd), .S(_433__bF_buf0) );
DFFSR DFFSR_105 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_430__5_), .Q(clgen_cnt_5_), .R(vdd), .S(_433__bF_buf3) );
DFFSR DFFSR_106 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf0), .D(_430__6_), .Q(clgen_cnt_6_), .R(vdd), .S(_433__bF_buf2) );
DFFSR DFFSR_107 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf0), .D(_430__7_), .Q(clgen_cnt_7_), .R(vdd), .S(_433__bF_buf1) );
DFFSR DFFSR_108 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf0), .D(_430__8_), .Q(clgen_cnt_8_), .R(vdd), .S(_433__bF_buf0) );
DFFSR DFFSR_109 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf0), .D(_430__9_), .Q(clgen_cnt_9_), .R(vdd), .S(_433__bF_buf3) );
DFFSR DFFSR_110 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf0), .D(_430__10_), .Q(clgen_cnt_10_), .R(vdd), .S(_433__bF_buf2) );
DFFSR DFFSR_111 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf0), .D(_430__11_), .Q(clgen_cnt_11_), .R(vdd), .S(_433__bF_buf1) );
DFFSR DFFSR_112 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf0), .D(_430__12_), .Q(clgen_cnt_12_), .R(vdd), .S(_433__bF_buf0) );
DFFSR DFFSR_113 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf0), .D(_430__13_), .Q(clgen_cnt_13_), .R(vdd), .S(_433__bF_buf3) );
DFFSR DFFSR_114 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf0), .D(_430__14_), .Q(clgen_cnt_14_), .R(vdd), .S(_433__bF_buf2) );
DFFSR DFFSR_115 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf0), .D(_430__15_), .Q(clgen_cnt_15_), .R(vdd), .S(_433__bF_buf1) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .Y(_1490_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .Y(_1491_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .Y(_1492_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1492_), .Y(_1493_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .B(_1493_), .Y(_1494_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1494_), .Y(_1495_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(shift_cnt_5_), .Y(_1496_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_6_), .B(_1496_), .Y(_1497_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .Y(_1498_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_7_), .B(_1498_), .Y(clgen_last_clk) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_423_), .Y(_1499_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(clgen_neg_edge), .B(clgen_pos_edge), .S(shift_tx_negedge), .Y(_1500_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(clgen_last_clk), .Y(_1501_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf2), .Y(_1502_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .Y(_1503_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .B(_1503_), .Y(_1504_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .Y(_1505_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf3), .B(char_len_0_), .C(_1503_), .Y(_1506_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1502__bF_buf2), .C(_1506_), .Y(_1507_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .Y(_1508_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1508_), .Y(_1509_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1510_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_1_), .B(char_len_1_), .Y(_1511_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(_1505_), .Y(_1512_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(char_len_0_), .C(_1511_), .Y(_1513_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .Y(_1514_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1512_), .C(lsb_bF_buf1), .Y(_1515_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf0), .B(_1510_), .C(_1515_), .Y(_1516_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .Y(_1517_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .C(shift_cnt_2_), .Y(_1518_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .B(_1493_), .Y(_1519_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .B(char_len_2_), .Y(_1520_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(char_len_1_), .Y(_1521_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_1_), .B(_1521_), .C(_1513_), .Y(_1522_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1522_), .Y(_1523_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .Y(_1524_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1522_), .Y(_1525_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1525_), .C(lsb_bF_buf3), .Y(_1526_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf2), .B(_1519_), .C(_1526_), .Y(_1527_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(char_len_2_), .Y(_1528_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .B(_1528_), .C(_1523_), .Y(_1529_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .B(char_len_3_), .Y(_1530_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1530_), .Y(_1531_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1532_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .Y(_1533_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .B(shift_cnt_2_), .C(shift_cnt_3_), .Y(_1534_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1534_), .Y(_1535_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf1), .B(_1535_), .Y(_1536_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1502__bF_buf0), .C(_1536_), .Y(_1537_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .Y(_1538_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_6_), .Y(_1539_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1539_), .Y(_1540_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .Y(_1541_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_5_), .B(_1541_), .Y(_1542_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .Y(_1543_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(_1543_), .Y(_1544_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_5_), .Y(_1545_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .B(_1545_), .Y(_1546_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1546_), .Y(_1547_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1547_), .C(_1542_), .Y(_1548_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .B(_1490_), .Y(_1549_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1549_), .Y(_1550_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(char_len_3_), .Y(_1551_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .Y(_1552_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1552_), .B(char_len_3_), .C(_1529_), .Y(_1553_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .B(_1551_), .C(_1553_), .Y(_1554_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1547_), .C(_1554_), .Y(_1555_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1555_), .Y(_1556_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_6_), .B(char_len_6_), .Y(_1557_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .B(_1556_), .Y(_1558_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .Y(_1559_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1555_), .C(_1559_), .Y(_1560_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1560_), .C(lsb_bF_buf1), .Y(_1561_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf0), .B(_1540_), .C(_1561__bF_buf6), .Y(_1562_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1554_), .Y(_1563_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(_1543_), .C(_1563_), .Y(_1564_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1547_), .Y(_1565_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(shift_cnt_4_), .C(shift_cnt_5_), .Y(_1566_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1496_), .Y(_1567_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf3), .B(_1567_), .Y(_1568_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1502__bF_buf2), .C(_1568_), .Y(_1569_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(rx_43_), .Y(_1570_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(rx_59_), .Y(_1571_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1550_), .Y(_1572_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(shift_cnt_3_), .C(shift_cnt_4_), .Y(_1573_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1573_), .Y(_1574_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf1), .B(_1574_), .Y(_1575_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_1502__bF_buf0), .C(_1575_), .Y(_1576_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1571_), .S(_1576__bF_buf4), .Y(_1577_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1569__bF_buf4), .Y(_1578_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1547_), .Y(_1579_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .Y(_1580_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf3), .B(_1580_), .Y(_1581_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1502__bF_buf2), .C(_1581_), .Y(_1582_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(rx_11_), .Y(_1583_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(rx_27_), .Y(_1584_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .B(_1584_), .S(_1576__bF_buf3), .Y(_1585_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1582__bF_buf4), .Y(_1586_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1578_), .B(_1586_), .C(_1562_), .Y(_1587_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1588_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(rx_107_), .Y(_1589_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(rx_123_), .Y(_1590_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(_1590_), .S(_1576__bF_buf2), .Y(_1591_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1591_), .B(_1569__bF_buf3), .Y(_1592_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(rx_75_), .Y(_1593_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(rx_91_), .Y(_1594_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1594_), .S(_1576__bF_buf1), .Y(_1595_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .B(_1582__bF_buf3), .Y(_1596_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .B(_1596_), .C(_1588_), .Y(_1597_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1587_), .C(_1538_), .Y(_1598_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(rx_115_), .Y(_1599_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf1), .B(_1540_), .Y(_1600_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1555_), .C(_1557_), .Y(_1601_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1556_), .Y(_1602_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1601_), .C(lsb_bF_buf3), .Y(_1603_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1604_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(rx_51_), .Y(_1605_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1540_), .B(lsb_bF_buf2), .Y(_1606_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .B(_1606__bF_buf5), .C(_1561__bF_buf5), .Y(_1607_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1604_), .C(_1607_), .Y(_1608_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(rx_19_), .Y(_1609_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1606__bF_buf4), .C(_1561__bF_buf4), .Y(_1610_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(rx_83_), .Y(_1611_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1612_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1610_), .C(_1612_), .Y(_1613_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1613_), .C(_1576__bF_buf0), .Y(_1614_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(_1576__bF_buf4), .Y(_1615_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(rx_3_), .Y(_1616_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1606__bF_buf3), .C(_1561__bF_buf3), .Y(_1617_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(rx_67_), .Y(_1618_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1619_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1617_), .C(_1619_), .Y(_1620_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(rx_99_), .Y(_1621_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1622_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(rx_35_), .Y(_1623_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1606__bF_buf2), .C(_1561__bF_buf2), .Y(_1624_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf1), .B(_1622_), .C(_1624_), .Y(_1625_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_1625_), .C(_1615_), .Y(_1626_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1626_), .C(_1537_), .Y(_1627_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1598_), .C(_1627_), .Y(_1628_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .Y(_1629_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(rx_31_), .Y(_1630_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1630_), .B(_1606__bF_buf1), .C(_1561__bF_buf1), .Y(_1631_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(rx_95_), .Y(_1632_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1633_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1633_), .C(_1569__bF_buf0), .Y(_1634_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(rx_127_), .Y(_1635_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1636_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(rx_63_), .Y(_1637_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1606__bF_buf0), .C(_1561__bF_buf0), .Y(_1638_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1638_), .C(_1582__bF_buf0), .Y(_1639_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1639_), .C(_1615_), .Y(_1640_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(rx_15_), .Y(_1641_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(_1606__bF_buf5), .C(_1561__bF_buf6), .Y(_1642_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(rx_79_), .Y(_1643_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1644_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1642_), .B(_1644_), .C(_1569__bF_buf4), .Y(_1645_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(rx_47_), .Y(_1646_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1606__bF_buf4), .C(_1561__bF_buf5), .Y(_1647_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(rx_111_), .Y(_1648_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1649_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_1649_), .C(_1582__bF_buf4), .Y(_1650_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .B(_1650_), .C(_1576__bF_buf3), .Y(_1651_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1640_), .C(_1651_), .Y(_1652_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(rx_119_), .Y(_1653_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1654_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(rx_55_), .Y(_1655_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1606__bF_buf3), .C(_1561__bF_buf4), .Y(_1656_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf3), .B(_1654_), .C(_1656_), .Y(_1657_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(rx_23_), .Y(_1658_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1658_), .B(_1606__bF_buf2), .C(_1561__bF_buf3), .Y(_1659_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(rx_87_), .Y(_1660_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1661_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf3), .B(_1659_), .C(_1661_), .Y(_1662_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1662_), .C(_1576__bF_buf2), .Y(_1663_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(rx_103_), .Y(_1664_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1665_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(rx_39_), .Y(_1666_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1606__bF_buf1), .C(_1561__bF_buf2), .Y(_1667_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1665_), .C(_1667_), .Y(_1668_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(rx_7_), .Y(_1669_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1606__bF_buf0), .C(_1561__bF_buf1), .Y(_1670_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(rx_71_), .Y(_1671_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1672_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1670_), .C(_1672_), .Y(_1673_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1673_), .C(_1615_), .Y(_1674_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(_1674_), .C(_1537_), .Y(_1675_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1652_), .C(_1675_), .Y(_1676_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .B(_1628_), .C(_1676_), .Y(_1677_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(rx_9_), .Y(_1678_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .B(_1576__bF_buf1), .Y(_1679_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(rx_25_), .B(_1576__bF_buf0), .C(_1679_), .Y(_1680_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1680_), .Y(_1681_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(rx_41_), .Y(_1682_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(rx_57_), .Y(_1683_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(_1683_), .S(_1576__bF_buf4), .Y(_1684_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1684_), .B(_1582__bF_buf0), .Y(_1685_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_1685_), .C(_1588_), .Y(_1686_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(rx_73_), .Y(_1687_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(rx_89_), .Y(_1688_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1688_), .S(_1576__bF_buf3), .Y(_1689_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1569__bF_buf1), .Y(_1690_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(rx_105_), .Y(_1691_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(rx_121_), .Y(_1692_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(_1692_), .S(_1576__bF_buf2), .Y(_1693_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_1582__bF_buf4), .Y(_1694_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .B(_1690_), .C(_1562_), .Y(_1695_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1686_), .C(_1629_), .Y(_1696_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(rx_109_), .Y(_1697_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(rx_125_), .Y(_1698_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1698_), .S(_1576__bF_buf1), .Y(_1699_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .B(_1569__bF_buf0), .Y(_1700_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(rx_77_), .Y(_1701_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(rx_93_), .Y(_1702_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_1702_), .S(_1576__bF_buf0), .Y(_1703_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_1582__bF_buf3), .Y(_1704_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1700_), .B(_1704_), .C(_1588_), .Y(_1705_) );
INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(rx_45_), .Y(_1706_) );
INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(rx_61_), .Y(_1707_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1707_), .S(_1576__bF_buf4), .Y(_1708_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1708_), .B(_1569__bF_buf4), .Y(_1709_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(rx_13_), .Y(_1710_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(rx_29_), .Y(_1711_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1710_), .B(_1711_), .S(_1576__bF_buf3), .Y(_1712_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1712_), .B(_1582__bF_buf2), .Y(_1713_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(_1713_), .C(_1562_), .Y(_1714_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1527_), .C(_1705_), .Y(_1715_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1696_), .B(_1715_), .C(_1538_), .Y(_1716_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(rx_17_), .Y(_1717_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(_1606__bF_buf5), .C(_1561__bF_buf0), .Y(_1718_) );
INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(rx_81_), .Y(_1719_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1720_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1718_), .C(_1720_), .Y(_1721_) );
INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(rx_113_), .Y(_1722_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1723_) );
INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(rx_49_), .Y(_1724_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_1606__bF_buf4), .C(_1561__bF_buf6), .Y(_1725_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf3), .B(_1723_), .C(_1725_), .Y(_1726_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1721_), .C(_1726_), .Y(_1727_) );
INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(rx_97_), .Y(_1728_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1729_) );
INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(rx_33_), .Y(_1730_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1606__bF_buf3), .C(_1561__bF_buf5), .Y(_1731_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1729_), .C(_1731_), .Y(_1732_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(rx_1_), .Y(_1733_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1606__bF_buf2), .C(_1561__bF_buf4), .Y(_1734_) );
INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(rx_65_), .Y(_1735_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1736_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf0), .B(_1734_), .C(_1736_), .Y(_1737_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1576__bF_buf2), .B(_1732_), .C(_1737_), .Y(_1738_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1727_), .C(_1738_), .Y(_1739_) );
INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(rx_117_), .Y(_1740_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1741_) );
INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(rx_53_), .Y(_1742_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(_1606__bF_buf1), .C(_1561__bF_buf3), .Y(_1743_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf1), .B(_1741_), .C(_1743_), .Y(_1744_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(rx_21_), .Y(_1745_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(_1606__bF_buf0), .C(_1561__bF_buf2), .Y(_1746_) );
INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(rx_85_), .Y(_1747_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1748_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf4), .B(_1746_), .C(_1748_), .Y(_1749_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1744_), .C(_1749_), .Y(_1750_) );
INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(rx_101_), .Y(_1751_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1752_) );
INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(rx_37_), .Y(_1753_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1606__bF_buf5), .C(_1561__bF_buf1), .Y(_1754_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf0), .B(_1752_), .C(_1754_), .Y(_1755_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(rx_5_), .Y(_1756_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .B(_1606__bF_buf4), .C(_1561__bF_buf0), .Y(_1757_) );
INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(rx_69_), .Y(_1758_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1759_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf3), .B(_1757_), .C(_1759_), .Y(_1760_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1576__bF_buf1), .B(_1755_), .C(_1760_), .Y(_1761_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1750_), .C(_1761_), .Y(_1762_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1739_), .C(_1762_), .Y(_1763_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1716_), .C(_1763_), .Y(_1764_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1764_), .C(_1677_), .Y(_1765_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1766_) );
INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(rx_126_), .Y(_1767_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1768_) );
INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(rx_62_), .Y(_1769_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(_1606__bF_buf3), .C(_1561__bF_buf6), .Y(_1770_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf4), .B(_1768_), .C(_1770_), .Y(_1771_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(rx_30_), .Y(_1772_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1772_), .B(_1606__bF_buf2), .C(_1561__bF_buf5), .Y(_1773_) );
INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(rx_94_), .Y(_1774_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1775_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1773_), .C(_1775_), .Y(_1776_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_1776_), .C(_1576__bF_buf0), .Y(_1777_) );
INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(rx_110_), .Y(_1778_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1779_) );
INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(rx_46_), .Y(_1780_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1606__bF_buf1), .C(_1561__bF_buf4), .Y(_1781_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf3), .B(_1779_), .C(_1781_), .Y(_1782_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(rx_14_), .Y(_1783_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1606__bF_buf0), .C(_1561__bF_buf3), .Y(_1784_) );
INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(rx_78_), .Y(_1785_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1786_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1784_), .C(_1786_), .Y(_1787_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1782_), .B(_1787_), .C(_1615_), .Y(_1788_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_1788_), .C(_1538_), .Y(_1789_) );
INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(rx_118_), .Y(_1790_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1791_) );
INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(rx_54_), .Y(_1792_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1606__bF_buf5), .C(_1561__bF_buf2), .Y(_1793_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1791_), .C(_1793_), .Y(_1794_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(rx_22_), .Y(_1795_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(_1606__bF_buf4), .C(_1561__bF_buf1), .Y(_1796_) );
INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(rx_86_), .Y(_1797_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1798_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf0), .B(_1796_), .C(_1798_), .Y(_1799_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_1799_), .C(_1576__bF_buf4), .Y(_1800_) );
INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(rx_102_), .Y(_1801_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1802_) );
INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(rx_38_), .Y(_1803_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1606__bF_buf3), .C(_1561__bF_buf0), .Y(_1804_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf1), .B(_1802_), .C(_1804_), .Y(_1805_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(rx_6_), .Y(_1806_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1806_), .B(_1606__bF_buf2), .C(_1561__bF_buf6), .Y(_1807_) );
INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(rx_70_), .Y(_1808_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1809_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf4), .B(_1807_), .C(_1809_), .Y(_1810_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_1810_), .C(_1615_), .Y(_1811_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1811_), .C(_1537_), .Y(_1812_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1789_), .C(_1812_), .Y(_1813_) );
INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(rx_122_), .Y(_1814_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1815_) );
INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(rx_58_), .Y(_1816_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1606__bF_buf1), .C(_1561__bF_buf5), .Y(_1817_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf0), .B(_1815_), .C(_1817_), .Y(_1818_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(rx_26_), .Y(_1819_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(_1606__bF_buf0), .C(_1561__bF_buf4), .Y(_1820_) );
INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(rx_90_), .Y(_1821_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1822_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf3), .B(_1820_), .C(_1822_), .Y(_1823_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1823_), .C(_1576__bF_buf3), .Y(_1824_) );
INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(rx_106_), .Y(_1825_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1826_) );
INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(rx_42_), .Y(_1827_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1606__bF_buf5), .C(_1561__bF_buf3), .Y(_1828_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf4), .B(_1826_), .C(_1828_), .Y(_1829_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(rx_10_), .Y(_1830_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(_1606__bF_buf4), .C(_1561__bF_buf2), .Y(_1831_) );
INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(rx_74_), .Y(_1832_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1833_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1831_), .C(_1833_), .Y(_1834_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(_1834_), .C(_1615_), .Y(_1835_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1824_), .B(_1835_), .C(_1538_), .Y(_1836_) );
INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(rx_114_), .Y(_1837_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1838_) );
INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(rx_50_), .Y(_1839_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1606__bF_buf3), .C(_1561__bF_buf1), .Y(_1840_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf3), .B(_1838_), .C(_1840_), .Y(_1841_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(rx_18_), .Y(_1842_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1606__bF_buf2), .C(_1561__bF_buf0), .Y(_1843_) );
INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(rx_82_), .Y(_1844_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1845_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1843_), .C(_1845_), .Y(_1846_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(_1846_), .C(_1576__bF_buf2), .Y(_1847_) );
INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(rx_98_), .Y(_1848_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1849_) );
INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(rx_34_), .Y(_1850_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1606__bF_buf1), .C(_1561__bF_buf6), .Y(_1851_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1849_), .C(_1851_), .Y(_1852_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(rx_2_), .Y(_1853_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1606__bF_buf0), .C(_1561__bF_buf5), .Y(_1854_) );
INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(rx_66_), .Y(_1855_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1856_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf0), .B(_1854_), .C(_1856_), .Y(_1857_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1857_), .C(_1615_), .Y(_1858_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(_1858_), .C(_1537_), .Y(_1859_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1836_), .C(_1859_), .Y(_1860_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .B(_1813_), .C(_1860_), .Y(_1861_) );
INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(rx_108_), .Y(_1862_) );
INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(rx_124_), .Y(_1863_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1863_), .S(_1576__bF_buf1), .Y(_1864_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1569__bF_buf1), .Y(_1865_) );
INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(rx_76_), .Y(_1866_) );
INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(rx_92_), .Y(_1867_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_1867_), .S(_1576__bF_buf0), .Y(_1868_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1582__bF_buf4), .Y(_1869_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1865_), .C(_1869_), .Y(_1870_) );
INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(rx_44_), .Y(_1871_) );
INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(rx_60_), .Y(_1872_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1871_), .B(_1872_), .S(_1576__bF_buf4), .Y(_1873_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1873_), .B(_1569__bF_buf0), .Y(_1874_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(rx_12_), .Y(_1875_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(rx_28_), .Y(_1876_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1876_), .S(_1576__bF_buf3), .Y(_1877_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1877_), .B(_1582__bF_buf3), .Y(_1878_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1874_), .B(_1878_), .C(_1588_), .Y(_1879_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1870_), .C(_1879_), .Y(_1880_) );
INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(rx_100_), .Y(_1881_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1882_) );
INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(rx_36_), .Y(_1883_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(_1606__bF_buf5), .C(_1561__bF_buf4), .Y(_1884_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf4), .B(_1882_), .C(_1884_), .Y(_1885_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(rx_4_), .Y(_1886_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(_1606__bF_buf4), .C(_1561__bF_buf3), .Y(_1887_) );
INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(rx_68_), .Y(_1888_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1889_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1887_), .C(_1889_), .Y(_1890_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_1890_), .C(_1615_), .Y(_1891_) );
INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(rx_116_), .Y(_1892_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1893_) );
INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(rx_52_), .Y(_1894_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1606__bF_buf3), .C(_1561__bF_buf2), .Y(_1895_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf3), .B(_1893_), .C(_1895_), .Y(_1896_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(rx_20_), .Y(_1897_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_1606__bF_buf2), .C(_1561__bF_buf1), .Y(_1898_) );
INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(rx_84_), .Y(_1899_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1900_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf1), .B(_1898_), .C(_1900_), .Y(_1901_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_1901_), .C(_1576__bF_buf2), .Y(_1902_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1902_), .C(_1537_), .Y(_1903_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .B(_1903_), .C(_1527_), .Y(_1904_) );
INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(rx_120_), .Y(_1905_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1906_) );
INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(rx_56_), .Y(_1907_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_1606__bF_buf1), .C(_1561__bF_buf0), .Y(_1908_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf2), .B(_1906_), .C(_1908_), .Y(_1909_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(rx_24_), .Y(_1910_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_1606__bF_buf0), .C(_1561__bF_buf6), .Y(_1911_) );
INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(rx_88_), .Y(_1912_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1913_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf0), .B(_1911_), .C(_1913_), .Y(_1914_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1909_), .B(_1914_), .C(_1576__bF_buf1), .Y(_1915_) );
INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(rx_104_), .Y(_1916_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1600__bF_buf5), .C(_1603__bF_buf5), .Y(_1917_) );
INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(rx_40_), .Y(_1918_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(_1606__bF_buf5), .C(_1561__bF_buf5), .Y(_1919_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf1), .B(_1917_), .C(_1919_), .Y(_1920_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(rx_8_), .Y(_1921_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_1606__bF_buf4), .C(_1561__bF_buf4), .Y(_1922_) );
INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(rx_72_), .Y(_1923_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_1600__bF_buf4), .C(_1603__bF_buf4), .Y(_1924_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf4), .B(_1922_), .C(_1924_), .Y(_1925_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1925_), .C(_1615_), .Y(_1926_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_1926_), .C(_1538_), .Y(_1927_) );
INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(rx_112_), .Y(_1928_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_1600__bF_buf3), .C(_1603__bF_buf3), .Y(_1929_) );
INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(rx_48_), .Y(_1930_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1606__bF_buf3), .C(_1561__bF_buf3), .Y(_1931_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf0), .B(_1929_), .C(_1931_), .Y(_1932_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(rx_16_), .Y(_1933_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_1606__bF_buf2), .C(_1561__bF_buf2), .Y(_1934_) );
INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(rx_80_), .Y(_1935_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_1600__bF_buf2), .C(_1603__bF_buf2), .Y(_1936_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf3), .B(_1934_), .C(_1936_), .Y(_1937_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1937_), .C(_1576__bF_buf0), .Y(_1938_) );
INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(rx_96_), .Y(_1939_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .B(_1600__bF_buf1), .C(_1603__bF_buf1), .Y(_1940_) );
INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(rx_32_), .Y(_1941_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1606__bF_buf1), .C(_1561__bF_buf1), .Y(_1942_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1569__bF_buf4), .B(_1940_), .C(_1942_), .Y(_1943_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(rx_0_), .Y(_1944_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(_1606__bF_buf0), .C(_1561__bF_buf0), .Y(_1945_) );
INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(rx_64_), .Y(_1946_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1600__bF_buf0), .C(_1603__bF_buf0), .Y(_1947_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1582__bF_buf2), .B(_1945_), .C(_1947_), .Y(_1948_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1948_), .C(_1615_), .Y(_1949_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1949_), .C(_1537_), .Y(_1950_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1927_), .B(_1950_), .C(_1629_), .Y(_1951_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1951_), .B(_1904_), .C(_1516_), .Y(_1952_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1766_), .B(_1861_), .C(_1952_), .Y(_1953_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1765_), .C(_1953_), .Y(_1954_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .B(_1501_), .C(_1954_), .Y(_545_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .Y(_1955_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1540_), .Y(_1956_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .B(_1539_), .C(lsb_bF_buf1), .Y(_1957_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .C(rx_negedge), .Y(_1958_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .Y(_1959_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .B(shift_cnt_3_), .C(_1959_), .Y(_1960_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1491_), .C(_1552_), .Y(_1961_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1961_), .C(_1960_), .Y(_1962_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(shift_cnt_1_), .Y(_1963_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1955_), .C(shift_cnt_2_), .Y(_1964_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .B(_1491_), .Y(_1965_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1965_), .C(_1964_), .Y(_1966_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1966_), .Y(_1967_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(_1960_), .C(_1551_), .Y(_1968_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1962_), .C(_1968_), .Y(_1969_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .B(_1963_), .C(_1533_), .Y(_1970_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_1_), .B(_1955_), .Y(_1971_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(char_len_1_), .B(_1971_), .C(_1970_), .Y(_1972_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(rx_negedge), .Y(_1973_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .B(_1973_), .Y(_1974_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1970_), .C(char_len_1_), .Y(_1975_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1975_), .B(_1974_), .C(_1972_), .Y(_1976_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .B(char_len_2_), .Y(_1977_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(char_len_3_), .B(_1961_), .C(_1960_), .Y(_1978_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1491_), .C(shift_cnt_3_), .Y(_1979_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .B(_1552_), .C(_1959_), .Y(_1980_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1979_), .C(_1980_), .Y(_1981_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1981_), .Y(_1982_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_1977_), .C(_1982_), .Y(_1983_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1983_), .Y(_1984_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1552_), .C(_1958_), .Y(_1985_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(shift_cnt_5_), .C(_1985_), .Y(_1986_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(_1985_), .C(shift_cnt_5_), .Y(_1987_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_1987_), .Y(_1988_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1988_), .C(_1541_), .Y(_1989_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .Y(_1990_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .B(_1987_), .C(_1990_), .Y(_1991_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1491_), .Y(_1992_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_1552_), .C(shift_cnt_4_), .Y(_1993_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1985_), .Y(_1994_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .B(_1994_), .C(_1993_), .Y(_1995_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(_1985_), .Y(_1996_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_1552_), .C(_1490_), .Y(_1997_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(_1996_), .C(_1997_), .Y(_1998_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1998_), .Y(_1999_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1989_), .C(_1999_), .Y(_2000_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1987_), .C(char_len_5_), .Y(_2001_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1995_), .C(_2001_), .Y(_2002_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1984_), .B(_2000_), .C(_2002_), .Y(_2003_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1557_), .Y(_2004_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_2003_), .Y(_2005_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_1_), .Y(_2006_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_1955_), .Y(_2007_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1492_), .C(rx_negedge), .Y(_2008_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .B(_2008_), .C(_1521_), .Y(_2009_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .B(char_len_0_), .Y(_2010_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_2007_), .C(_2008_), .Y(_2011_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(_2011_), .C(_2009_), .Y(_2012_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .B(_1528_), .Y(_2013_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1968_), .Y(_2014_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2013_), .C(_2014_), .Y(_2015_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(_2015_), .Y(_2016_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1986_), .C(_1988_), .Y(_2017_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1998_), .Y(_2018_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_2001_), .C(_2018_), .Y(_2019_) );
INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .Y(_2020_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_2017_), .C(_1989_), .Y(_2021_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_2016_), .C(_2021_), .Y(_2022_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .Y(_2023_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2023_), .B(_2022_), .C(_1502__bF_buf0), .Y(_2024_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1957_), .C(_2024_), .D(_2005_), .Y(_2025_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1955_), .C(_1502__bF_buf3), .Y(_2026_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1567_), .C(_2026_), .Y(_2027_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_2001_), .B(_2017_), .Y(_2028_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .Y(_2029_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1983_), .C(_1999_), .Y(_2030_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(_2020_), .C(_2029_), .Y(_2031_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(_2018_), .C(_2015_), .Y(_2032_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_1995_), .C(_2032_), .Y(_2033_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2031_), .C(_1502__bF_buf2), .Y(_2034_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1574_), .Y(_2035_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(_1955_), .C(_2035_), .Y(_2036_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(lsb_bF_buf0), .Y(_2037_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1999_), .C(_1983_), .Y(_2038_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf3), .B(_2038_), .C(_2032_), .Y(_2039_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2037_), .Y(_2040_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2027_), .C(_2034_), .Y(_2041_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_2041__bF_buf3), .Y(_2042_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2025__bF_buf7), .B(_2042_), .Y(_2043_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .B(rx_negedge), .C(lsb_bF_buf2), .Y(_2044_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(rx_negedge), .C(_2044_), .Y(_2045_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .Y(_2046_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_1977_), .Y(_2047_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1966_), .C(_2047_), .Y(_2048_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_2048_), .C(_1502__bF_buf1), .Y(_2049_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_2048_), .C(_2049_), .Y(_2050_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2050_), .Y(_2051_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1977_), .B(_2012_), .Y(_2052_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1519_), .B(rx_negedge), .C(_1965_), .Y(_2053_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf0), .B(_2053_), .Y(_2054_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(_1502__bF_buf3), .C(_2054_), .Y(_2055_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2051_), .Y(_2056_) );
INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .Y(_2057_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1492_), .C(_1955_), .Y(_2058_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_1955_), .C(_2058_), .Y(_2059_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1502__bF_buf2), .B(_2059_), .Y(_2060_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_2011_), .B(_1972_), .Y(_2061_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_2061_), .B(_2010_), .Y(_2062_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf1), .B(_2062_), .Y(_2063_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2063_), .Y(_2064_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2065_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .B(_1502__bF_buf1), .Y(_2066_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .B(_2066_), .Y(_2067_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_2067_), .Y(_2068_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2065_), .Y(_2069_) );
INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(_2069_), .Y(_2070_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2057_), .Y(_2071_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2043_), .Y(_2072_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2051_), .Y(_2073_) );
INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(_2073_), .Y(_2074_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1957_), .B(_1956_), .Y(_2075_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2023_), .B(_2022_), .Y(_2076_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2003_), .B(_2004_), .C(lsb_bF_buf0), .Y(_2077_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_2076_), .C(_2075_), .Y(_2078_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(rx_33_), .B(_2078__bF_buf7), .Y(_2079_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf3), .B(_2036_), .C(_2039_), .Y(_2080_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .B(_2080_), .C(_2034_), .Y(_2081_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(rx_97_), .B(_2025__bF_buf6), .C(_2081__bF_buf3), .Y(_2082_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(rx_49_), .B(_2078__bF_buf6), .Y(_2083_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(rx_113_), .B(_2025__bF_buf5), .C(_2041__bF_buf2), .Y(_2084_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2079_), .C(_2083_), .D(_2084_), .Y(_2085_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(rx_65_), .B(_2025__bF_buf4), .Y(_2086_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .Y(_2087_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(_2020_), .C(_2028_), .Y(_2088_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2029_), .B(_1995_), .C(_2032_), .Y(_2089_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf2), .B(_2089_), .C(_2088_), .Y(_2090_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_2090_), .C(_2080_), .Y(_2091_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_1_), .C(_2091__bF_buf3), .Y(_2092_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(rx_81_), .B(_2025__bF_buf3), .Y(_2093_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_2090_), .C(_2040_), .Y(_2094_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_17_), .C(_2094__bF_buf3), .Y(_2095_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_2086_), .C(_2093_), .D(_2095_), .Y(_2096_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2085_), .B(_2096_), .C(_2074_), .Y(_2097_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(rx_45_), .B(_2078__bF_buf3), .Y(_2098_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(rx_109_), .B(_2025__bF_buf2), .C(_2081__bF_buf2), .Y(_2099_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(rx_61_), .B(_2078__bF_buf2), .Y(_2100_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(rx_125_), .B(_2025__bF_buf1), .C(_2041__bF_buf1), .Y(_2101_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2098_), .C(_2100_), .D(_2101_), .Y(_2102_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(rx_77_), .B(_2025__bF_buf0), .Y(_2103_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_13_), .C(_2091__bF_buf2), .Y(_2104_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(rx_93_), .B(_2025__bF_buf7), .Y(_2105_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_29_), .C(_2094__bF_buf2), .Y(_2106_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2104_), .B(_2103_), .C(_2105_), .D(_2106_), .Y(_2107_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2102_), .B(_2107_), .C(_2056_), .Y(_2108_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(_2108_), .Y(_2109_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .Y(_2110_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2110_), .Y(_2111_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(rx_37_), .B(_2078__bF_buf7), .Y(_2112_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(rx_101_), .B(_2025__bF_buf6), .C(_2081__bF_buf1), .Y(_2113_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(rx_53_), .B(_2078__bF_buf6), .Y(_2114_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(rx_117_), .B(_2025__bF_buf5), .C(_2041__bF_buf0), .Y(_2115_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2112_), .C(_2114_), .D(_2115_), .Y(_2116_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(rx_69_), .B(_2025__bF_buf4), .Y(_2117_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_5_), .C(_2091__bF_buf1), .Y(_2118_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(rx_85_), .B(_2025__bF_buf3), .Y(_2119_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_21_), .C(_2094__bF_buf1), .Y(_2120_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2117_), .C(_2119_), .D(_2120_), .Y(_2121_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2121_), .C(_2111_), .Y(_2122_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2110_), .Y(_2123_) );
INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .Y(_2124_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(rx_41_), .B(_2078__bF_buf3), .Y(_2125_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(rx_105_), .B(_2025__bF_buf2), .C(_2081__bF_buf0), .Y(_2126_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(rx_57_), .B(_2078__bF_buf2), .Y(_2127_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(rx_121_), .B(_2025__bF_buf1), .C(_2041__bF_buf3), .Y(_2128_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(_2125_), .C(_2127_), .D(_2128_), .Y(_2129_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(rx_73_), .B(_2025__bF_buf0), .Y(_2130_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_9_), .C(_2091__bF_buf0), .Y(_2131_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(rx_89_), .B(_2025__bF_buf7), .Y(_2132_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_25_), .C(_2094__bF_buf0), .Y(_2133_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2130_), .C(_2132_), .D(_2133_), .Y(_2134_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(_2134_), .C(_2124_), .Y(_2135_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_2122_), .B(_2135_), .Y(_2136_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2064_), .Y(_2137_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2136_), .C(_2137_), .Y(_2138_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(clgen_last_clk), .Y(_2139_) );
INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(clgen_pos_edge), .Y(_2140_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(clgen_neg_edge), .B(rx_negedge), .Y(_2141_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(rx_negedge), .C(_2141_), .Y(_2142_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(_424_), .C(_2142_), .Y(_2143_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(rx_32_), .B(_2078__bF_buf7), .Y(_2144_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(rx_96_), .B(_2025__bF_buf6), .C(_2081__bF_buf3), .Y(_2145_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(rx_48_), .B(_2078__bF_buf6), .Y(_2146_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(rx_112_), .B(_2025__bF_buf5), .C(_2041__bF_buf2), .Y(_2147_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(_2144_), .C(_2146_), .D(_2147_), .Y(_2148_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(rx_64_), .B(_2025__bF_buf4), .Y(_2149_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_0_), .C(_2091__bF_buf3), .Y(_2150_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(rx_80_), .B(_2025__bF_buf3), .Y(_2151_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_16_), .C(_2094__bF_buf3), .Y(_2152_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2149_), .C(_2151_), .D(_2152_), .Y(_548_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2148_), .B(_548_), .C(_2074_), .Y(_549_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(rx_44_), .B(_2078__bF_buf3), .Y(_550_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(rx_108_), .B(_2025__bF_buf2), .C(_2081__bF_buf2), .Y(_551_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(rx_60_), .B(_2078__bF_buf2), .Y(_552_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(rx_124_), .B(_2025__bF_buf1), .C(_2041__bF_buf1), .Y(_553_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_550_), .C(_552_), .D(_553_), .Y(_554_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(rx_76_), .B(_2025__bF_buf0), .Y(_555_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_12_), .C(_2091__bF_buf2), .Y(_556_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(rx_92_), .B(_2025__bF_buf7), .Y(_557_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_28_), .C(_2094__bF_buf2), .Y(_558_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_555_), .C(_557_), .D(_558_), .Y(_559_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_559_), .C(_2056_), .Y(_560_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_560_), .Y(_561_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(rx_36_), .B(_2078__bF_buf7), .Y(_562_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(rx_100_), .B(_2025__bF_buf6), .C(_2081__bF_buf1), .Y(_563_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(rx_52_), .B(_2078__bF_buf6), .Y(_564_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(rx_116_), .B(_2025__bF_buf5), .C(_2041__bF_buf0), .Y(_565_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_562_), .C(_564_), .D(_565_), .Y(_566_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(rx_68_), .B(_2025__bF_buf4), .Y(_567_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_4_), .C(_2091__bF_buf1), .Y(_568_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(rx_84_), .B(_2025__bF_buf3), .Y(_569_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_20_), .C(_2094__bF_buf1), .Y(_570_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_567_), .C(_569_), .D(_570_), .Y(_571_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_571_), .C(_2111_), .Y(_572_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(rx_40_), .B(_2078__bF_buf3), .Y(_573_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(rx_104_), .B(_2025__bF_buf2), .C(_2081__bF_buf0), .Y(_574_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(rx_56_), .B(_2078__bF_buf2), .Y(_575_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(rx_120_), .B(_2025__bF_buf1), .C(_2041__bF_buf3), .Y(_576_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_573_), .C(_575_), .D(_576_), .Y(_577_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(rx_72_), .B(_2025__bF_buf0), .Y(_578_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_8_), .C(_2091__bF_buf0), .Y(_579_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(rx_88_), .B(_2025__bF_buf7), .Y(_580_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_24_), .C(_2094__bF_buf0), .Y(_581_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_578_), .C(_580_), .D(_581_), .Y(_582_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_582_), .C(_2124_), .Y(_583_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_583_), .Y(_584_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_2067_), .B(_2064_), .Y(_585_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_584_), .C(_585_), .Y(_586_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2138_), .C(_586_), .Y(_587_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(rx_51_), .B(_2078__bF_buf7), .Y(_588_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(rx_115_), .B(_2025__bF_buf6), .C(_2041__bF_buf2), .Y(_589_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(rx_35_), .B(_2078__bF_buf6), .Y(_590_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(rx_99_), .B(_2025__bF_buf5), .C(_2081__bF_buf3), .Y(_591_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_590_), .C(_588_), .D(_589_), .Y(_592_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(rx_83_), .B(_2025__bF_buf4), .Y(_593_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_19_), .C(_2094__bF_buf3), .Y(_594_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(rx_67_), .B(_2025__bF_buf3), .Y(_595_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_3_), .C(_2091__bF_buf3), .Y(_596_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_593_), .C(_595_), .D(_596_), .Y(_597_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_597_), .C(_2074_), .Y(_598_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(rx_63_), .B(_2078__bF_buf3), .Y(_599_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(rx_127_), .B(_2025__bF_buf2), .C(_2041__bF_buf1), .Y(_600_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(rx_47_), .B(_2078__bF_buf2), .Y(_601_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(rx_111_), .B(_2025__bF_buf1), .C(_2081__bF_buf2), .Y(_602_) );
OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_601_), .C(_599_), .D(_600_), .Y(_603_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(rx_95_), .B(_2025__bF_buf0), .Y(_604_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_31_), .C(_2094__bF_buf2), .Y(_605_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(rx_79_), .B(_2025__bF_buf7), .Y(_606_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_15_), .C(_2091__bF_buf2), .Y(_607_) );
OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_604_), .C(_606_), .D(_607_), .Y(_608_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_608_), .C(_2056_), .Y(_609_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_609_), .Y(_610_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(rx_55_), .B(_2078__bF_buf7), .Y(_611_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(rx_119_), .B(_2025__bF_buf6), .C(_2041__bF_buf0), .Y(_612_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(rx_39_), .B(_2078__bF_buf6), .Y(_613_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(rx_103_), .B(_2025__bF_buf5), .C(_2081__bF_buf1), .Y(_614_) );
OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_613_), .C(_611_), .D(_612_), .Y(_615_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(rx_87_), .B(_2025__bF_buf4), .Y(_616_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_23_), .C(_2094__bF_buf1), .Y(_617_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(rx_71_), .B(_2025__bF_buf3), .Y(_618_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_7_), .C(_2091__bF_buf1), .Y(_619_) );
OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_616_), .C(_618_), .D(_619_), .Y(_620_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_620_), .C(_2111_), .Y(_621_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(rx_59_), .B(_2078__bF_buf3), .Y(_622_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(rx_123_), .B(_2025__bF_buf2), .C(_2041__bF_buf3), .Y(_623_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(rx_43_), .B(_2078__bF_buf2), .Y(_624_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(rx_107_), .B(_2025__bF_buf1), .C(_2081__bF_buf0), .Y(_625_) );
OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_624_), .C(_622_), .D(_623_), .Y(_626_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(rx_91_), .B(_2025__bF_buf0), .Y(_627_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_27_), .C(_2094__bF_buf0), .Y(_628_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(rx_75_), .B(_2025__bF_buf7), .Y(_629_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_11_), .C(_2091__bF_buf0), .Y(_630_) );
OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_627_), .C(_629_), .D(_630_), .Y(_631_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_631_), .C(_2124_), .Y(_632_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_632_), .Y(_633_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_633_), .C(_2069_), .Y(_634_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(rx_50_), .B(_2078__bF_buf7), .Y(_635_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(rx_114_), .B(_2025__bF_buf6), .C(_2041__bF_buf2), .Y(_636_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(rx_34_), .B(_2078__bF_buf6), .Y(_637_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(rx_98_), .B(_2025__bF_buf5), .C(_2081__bF_buf3), .Y(_638_) );
OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_637_), .C(_635_), .D(_636_), .Y(_639_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(rx_82_), .B(_2025__bF_buf4), .Y(_640_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_18_), .C(_2094__bF_buf3), .Y(_641_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(rx_66_), .B(_2025__bF_buf3), .Y(_642_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_2_), .C(_2091__bF_buf3), .Y(_643_) );
OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_640_), .C(_642_), .D(_643_), .Y(_644_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_644_), .C(_2074_), .Y(_645_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(rx_62_), .B(_2078__bF_buf3), .Y(_646_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(rx_126_), .B(_2025__bF_buf2), .C(_2041__bF_buf1), .Y(_647_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(rx_46_), .B(_2078__bF_buf2), .Y(_648_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(rx_110_), .B(_2025__bF_buf1), .C(_2081__bF_buf2), .Y(_649_) );
OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_648_), .C(_646_), .D(_647_), .Y(_650_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(rx_94_), .B(_2025__bF_buf0), .Y(_651_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_30_), .C(_2094__bF_buf2), .Y(_652_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(rx_78_), .B(_2025__bF_buf7), .Y(_653_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_14_), .C(_2091__bF_buf2), .Y(_654_) );
OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_651_), .C(_653_), .D(_654_), .Y(_655_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_655_), .C(_2056_), .Y(_656_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_656_), .Y(_657_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(rx_54_), .B(_2078__bF_buf7), .Y(_658_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(rx_118_), .B(_2025__bF_buf6), .C(_2041__bF_buf0), .Y(_659_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(rx_38_), .B(_2078__bF_buf6), .Y(_660_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(rx_102_), .B(_2025__bF_buf5), .C(_2081__bF_buf1), .Y(_661_) );
OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_660_), .C(_658_), .D(_659_), .Y(_662_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(rx_86_), .B(_2025__bF_buf4), .Y(_663_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(rx_22_), .C(_2094__bF_buf1), .Y(_664_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(rx_70_), .B(_2025__bF_buf3), .Y(_665_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(rx_6_), .C(_2091__bF_buf1), .Y(_666_) );
OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_663_), .C(_665_), .D(_666_), .Y(_667_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_667_), .C(_2111_), .Y(_668_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(rx_58_), .B(_2078__bF_buf3), .Y(_669_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(rx_122_), .B(_2025__bF_buf2), .C(_2041__bF_buf3), .Y(_670_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(rx_42_), .B(_2078__bF_buf2), .Y(_671_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(rx_106_), .B(_2025__bF_buf1), .C(_2081__bF_buf0), .Y(_672_) );
OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_671_), .C(_669_), .D(_670_), .Y(_673_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(rx_90_), .B(_2025__bF_buf0), .Y(_674_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf1), .B(rx_26_), .C(_2094__bF_buf0), .Y(_675_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(rx_74_), .B(_2025__bF_buf7), .Y(_676_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf0), .B(rx_10_), .C(_2091__bF_buf0), .Y(_677_) );
OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_674_), .C(_676_), .D(_677_), .Y(_678_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_678_), .C(_2124_), .Y(_679_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_679_), .Y(_680_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_2067_), .B(_2065_), .Y(_681_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_680_), .C(_681_), .Y(_682_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_682_), .Y(_683_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(miso_pad_i), .Y(_684_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_683_), .C(_684_), .Y(_685_) );
INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .Y(_686_) );
INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(shift_latch_3_), .Y(_687_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf2), .B(_687__bF_buf3), .Y(_688_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_2072_), .C(_688__bF_buf7), .Y(_689_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_2072_), .C(_689_), .Y(_690_) );
INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(shift_latch_2_), .Y(_691_) );
INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf1), .Y(_692_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(shift_latch_1_), .B(shift_latch_0_), .C(_692_), .Y(_693_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf0), .B(_691_), .C(_693__bF_buf5), .Y(_694_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[31]), .B(wb_sel_i_3_bF_buf4_), .Y(_695_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(wb_sel_i_3_bF_buf3_), .C(_695_), .Y(_696_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_696_), .C(_694__bF_buf7), .Y(_697_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_694__bF_buf6), .C(_690_), .D(_697_), .Y(_544__127_) );
INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(_681_), .Y(_698_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_2057_), .Y(_699_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2043_), .Y(_700_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(_700_), .C(_688__bF_buf5), .Y(_701_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf7), .B(_700_), .C(_701_), .Y(_702_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf2_), .B(wb_dat_i[30]), .Y(_703_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(wb_sel_i_3_bF_buf1_), .C(_703_), .Y(_704_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_704_), .C(_694__bF_buf5), .Y(_705_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(_694__bF_buf4), .C(_702_), .D(_705_), .Y(_544__126_) );
INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .Y(_706_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_2057_), .Y(_707_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_2043_), .Y(_708_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_708_), .C(_688__bF_buf3), .Y(_709_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_708_), .C(_709_), .Y(_710_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf0_), .B(wb_dat_i[29]), .Y(_711_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(wb_sel_i_3_bF_buf6_), .C(_711_), .Y(_712_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_712_), .C(_694__bF_buf3), .Y(_713_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_694__bF_buf2), .C(_710_), .D(_713_), .Y(_544__125_) );
INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_714_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_2057_), .Y(_715_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_2043_), .Y(_716_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_716_), .C(_688__bF_buf1), .Y(_717_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_716_), .C(_717_), .Y(_718_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf5_), .B(wb_dat_i[28]), .Y(_719_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(wb_sel_i_3_bF_buf4_), .C(_719_), .Y(_720_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_720_), .C(_694__bF_buf1), .Y(_721_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_694__bF_buf0), .C(_718_), .D(_721_), .Y(_544__124_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2123_), .Y(_722_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_2043_), .Y(_723_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_723_), .C(_688__bF_buf7), .Y(_724_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_723_), .C(_724_), .Y(_725_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf3_), .B(wb_dat_i[27]), .Y(_726_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(wb_sel_i_3_bF_buf2_), .C(_726_), .Y(_727_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_727_), .C(_694__bF_buf7), .Y(_728_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_694__bF_buf6), .C(_725_), .D(_728_), .Y(_544__123_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_2123_), .Y(_729_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_2043_), .Y(_730_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(_730_), .C(_688__bF_buf5), .Y(_731_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_730_), .C(_731_), .Y(_732_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf1_), .B(wb_dat_i[26]), .Y(_733_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(wb_sel_i_3_bF_buf0_), .C(_733_), .Y(_734_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_734_), .C(_694__bF_buf5), .Y(_735_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(_694__bF_buf4), .C(_732_), .D(_735_), .Y(_544__122_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_2123_), .Y(_736_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_2043_), .Y(_737_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_737_), .C(_688__bF_buf3), .Y(_738_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_737_), .C(_738_), .Y(_739_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf6_), .B(wb_dat_i[25]), .Y(_740_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(wb_sel_i_3_bF_buf5_), .C(_740_), .Y(_741_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_741_), .C(_694__bF_buf3), .Y(_742_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_694__bF_buf2), .C(_739_), .D(_742_), .Y(_544__121_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_2123_), .Y(_743_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_2043_), .Y(_744_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_744_), .C(_688__bF_buf1), .Y(_745_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf1), .B(_744_), .C(_745_), .Y(_746_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_3_bF_buf4_), .B(wb_dat_i[24]), .Y(_747_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(wb_sel_i_3_bF_buf3_), .C(_747_), .Y(_748_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_748_), .C(_694__bF_buf1), .Y(_749_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_694__bF_buf0), .C(_746_), .D(_749_), .Y(_544__120_) );
INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .Y(_750_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_750_), .Y(_751_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_751_), .Y(_752_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(_752_), .C(_688__bF_buf7), .Y(_753_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_752_), .C(_753_), .Y(_754_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[22]), .B(wb_sel_i_2_bF_buf4_), .Y(_755_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(wb_sel_i_2_bF_buf3_), .C(_755_), .Y(_756_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_756_), .C(_694__bF_buf7), .Y(_757_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(_694__bF_buf6), .C(_754_), .D(_757_), .Y(_544__118_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_750_), .Y(_758_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_758_), .Y(_759_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_759_), .C(_688__bF_buf5), .Y(_760_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_759_), .C(_760_), .Y(_761_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf2_), .B(wb_dat_i[21]), .Y(_762_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(wb_sel_i_2_bF_buf1_), .C(_762_), .Y(_763_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_763_), .C(_694__bF_buf5), .Y(_764_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_694__bF_buf4), .C(_761_), .D(_764_), .Y(_544__117_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_750_), .Y(_765_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_765_), .Y(_766_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_766_), .C(_688__bF_buf3), .Y(_767_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf7), .B(_766_), .C(_767_), .Y(_768_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf0_), .B(wb_dat_i[20]), .Y(_769_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(wb_sel_i_2_bF_buf6_), .C(_769_), .Y(_770_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_770_), .C(_694__bF_buf3), .Y(_771_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_694__bF_buf2), .C(_768_), .D(_771_), .Y(_544__116_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2073_), .Y(_772_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_2043_), .Y(_773_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_773_), .C(_688__bF_buf1), .Y(_774_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_773_), .C(_774_), .Y(_775_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf5_), .B(wb_dat_i[19]), .Y(_776_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(wb_sel_i_2_bF_buf4_), .C(_776_), .Y(_777_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_777_), .C(_694__bF_buf1), .Y(_778_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_694__bF_buf0), .C(_775_), .D(_778_), .Y(_544__115_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf3_), .B(wb_dat_i[18]), .Y(_779_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(wb_sel_i_2_bF_buf2_), .C(_779_), .Y(_780_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_688__bF_buf7), .Y(_781_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_2073_), .Y(_782_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_2043_), .Y(_783_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_783_), .Y(_784_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_685__bF_buf3), .Y(_785_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_783_), .C(_688__bF_buf6), .Y(_786_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_785_), .C(_781_), .Y(_787_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_691_), .Y(_788_) );
INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(_693__bF_buf4), .Y(_789_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf3), .B(_788__bF_buf4), .C(rx_114_), .Y(_790_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_694__bF_buf7), .C(_790_), .Y(_544__114_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_2073_), .Y(_791_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_2043_), .Y(_792_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(_792_), .C(_688__bF_buf5), .Y(_793_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_792_), .C(_793_), .Y(_794_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf1_), .B(wb_dat_i[17]), .Y(_795_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(wb_sel_i_2_bF_buf0_), .C(_795_), .Y(_796_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_796_), .C(_694__bF_buf6), .Y(_797_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(_694__bF_buf5), .C(_794_), .D(_797_), .Y(_544__113_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_2073_), .Y(_798_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_2043_), .Y(_799_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_799_), .C(_688__bF_buf3), .Y(_800_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_799_), .C(_800_), .Y(_801_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf6_), .B(wb_dat_i[16]), .Y(_802_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(wb_sel_i_2_bF_buf5_), .C(_802_), .Y(_803_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_803_), .C(_694__bF_buf4), .Y(_804_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_694__bF_buf3), .C(_801_), .D(_804_), .Y(_544__112_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[14]), .B(wb_sel_i_1_bF_buf1_), .Y(_805_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(wb_sel_i_1_bF_buf0_), .C(_805_), .Y(_806_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_688__bF_buf1), .Y(_807_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_2081__bF_buf3), .Y(_808_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2025__bF_buf6), .B(_808_), .Y(_809_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_809_), .Y(_810_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_699_), .Y(_811_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_810_), .Y(_812_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_685__bF_buf2), .Y(_813_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_812_), .Y(_814_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_814_), .C(_688__bF_buf0), .Y(_815_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_813_), .C(_807_), .Y(_816_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_788__bF_buf3), .C(rx_110_), .Y(_817_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_694__bF_buf2), .C(_817_), .Y(_544__110_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_809_), .Y(_818_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_818_), .C(_688__bF_buf7), .Y(_819_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_818_), .C(_819_), .Y(_820_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf7_), .B(wb_dat_i[13]), .Y(_821_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(wb_sel_i_1_bF_buf6_), .C(_821_), .Y(_822_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_822_), .C(_694__bF_buf1), .Y(_823_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_694__bF_buf0), .C(_820_), .D(_823_), .Y(_544__109_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_809_), .Y(_824_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_824_), .C(_688__bF_buf5), .Y(_825_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_824_), .C(_825_), .Y(_826_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf5_), .B(wb_dat_i[12]), .Y(_827_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(wb_sel_i_1_bF_buf4_), .C(_827_), .Y(_828_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_828_), .C(_694__bF_buf7), .Y(_829_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_694__bF_buf6), .C(_826_), .D(_829_), .Y(_544__108_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_809_), .Y(_830_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(_830_), .C(_688__bF_buf3), .Y(_831_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf1), .B(_830_), .C(_831_), .Y(_832_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf3_), .B(wb_dat_i[11]), .Y(_833_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(wb_sel_i_1_bF_buf2_), .C(_833_), .Y(_834_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_834_), .C(_694__bF_buf5), .Y(_835_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(_694__bF_buf4), .C(_832_), .D(_835_), .Y(_544__107_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf1_), .B(wb_dat_i[10]), .Y(_836_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(wb_sel_i_1_bF_buf0_), .C(_836_), .Y(_837_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_688__bF_buf1), .Y(_838_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_729_), .Y(_839_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_810_), .Y(_840_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_685__bF_buf1), .Y(_841_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_840_), .Y(_842_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(_842_), .C(_688__bF_buf0), .Y(_843_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_841_), .C(_838_), .Y(_844_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf1), .B(_788__bF_buf2), .C(rx_106_), .Y(_845_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_694__bF_buf3), .C(_845_), .Y(_544__106_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_809_), .Y(_846_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(_846_), .C(_688__bF_buf7), .Y(_847_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_846_), .C(_847_), .Y(_848_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf7_), .B(wb_dat_i[9]), .Y(_849_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(wb_sel_i_1_bF_buf6_), .C(_849_), .Y(_850_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_850_), .C(_694__bF_buf2), .Y(_851_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(_694__bF_buf1), .C(_848_), .D(_851_), .Y(_544__105_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_809_), .Y(_852_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_852_), .C(_688__bF_buf5), .Y(_853_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_852_), .C(_853_), .Y(_854_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf5_), .B(wb_dat_i[8]), .Y(_855_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(wb_sel_i_1_bF_buf4_), .C(_855_), .Y(_856_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_856_), .C(_694__bF_buf0), .Y(_857_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_694__bF_buf7), .C(_854_), .D(_857_), .Y(_544__104_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_751_), .Y(_858_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_858_), .C(_688__bF_buf3), .Y(_859_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf7), .B(_858_), .C(_859_), .Y(_860_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[6]), .B(wb_sel_i_0_bF_buf7_), .Y(_861_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(wb_sel_i_0_bF_buf6_), .C(_861_), .Y(_862_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_862_), .C(_694__bF_buf6), .Y(_863_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_694__bF_buf5), .C(_860_), .D(_863_), .Y(_544__102_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_758_), .Y(_864_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_864_), .C(_688__bF_buf1), .Y(_865_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_864_), .C(_865_), .Y(_866_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf5_), .B(wb_dat_i[5]), .Y(_867_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(wb_sel_i_0_bF_buf4_), .C(_867_), .Y(_868_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_868_), .C(_694__bF_buf4), .Y(_869_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_694__bF_buf3), .C(_866_), .D(_869_), .Y(_544__101_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_765_), .Y(_870_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(_870_), .C(_688__bF_buf7), .Y(_871_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_870_), .C(_871_), .Y(_872_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf3_), .B(wb_dat_i[4]), .Y(_873_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(wb_sel_i_0_bF_buf2_), .C(_873_), .Y(_874_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_874_), .C(_694__bF_buf2), .Y(_875_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(_694__bF_buf1), .C(_872_), .D(_875_), .Y(_544__100_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_809_), .Y(_876_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_876_), .C(_688__bF_buf5), .Y(_877_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_876_), .C(_877_), .Y(_878_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf1_), .B(wb_dat_i[3]), .Y(_879_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(wb_sel_i_0_bF_buf0_), .C(_879_), .Y(_880_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_880_), .C(_694__bF_buf0), .Y(_881_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_694__bF_buf7), .C(_878_), .D(_881_), .Y(_544__99_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_809_), .Y(_882_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_882_), .C(_688__bF_buf3), .Y(_883_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_882_), .C(_883_), .Y(_884_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf7_), .B(wb_dat_i[2]), .Y(_885_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(wb_sel_i_0_bF_buf6_), .C(_885_), .Y(_886_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_886_), .C(_694__bF_buf6), .Y(_887_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_694__bF_buf5), .C(_884_), .D(_887_), .Y(_544__98_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_809_), .Y(_888_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .B(_888_), .C(_688__bF_buf1), .Y(_889_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_888_), .C(_889_), .Y(_890_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf5_), .B(wb_dat_i[1]), .Y(_891_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .B(wb_sel_i_0_bF_buf4_), .C(_891_), .Y(_892_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_892_), .C(_694__bF_buf4), .Y(_893_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .B(_694__bF_buf3), .C(_890_), .D(_893_), .Y(_544__97_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_809_), .Y(_894_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .B(_894_), .C(_688__bF_buf7), .Y(_895_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf1), .B(_894_), .C(_895_), .Y(_896_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf3_), .B(wb_dat_i[0]), .Y(_897_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .B(wb_sel_i_0_bF_buf2_), .C(_897_), .Y(_898_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf6), .B(_898_), .C(_694__bF_buf2), .Y(_899_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .B(_694__bF_buf1), .C(_896_), .D(_899_), .Y(_544__96_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_2094__bF_buf3), .Y(_900_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_2025__bF_buf5), .B(_900_), .Y(_901_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf2), .B(clgen_enable_bF_buf8), .C(_699_), .Y(_902_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_903_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_903_), .Y(_904_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_904_), .C(_788__bF_buf1), .Y(_905_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_904_), .C(_905_), .Y(_906_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(wb_sel_i_3_bF_buf2_), .C(_703_), .Y(_907_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf0), .B(_907_), .C(_694__bF_buf0), .Y(_908_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_789__bF_buf3), .C(_906_), .D(_908_), .Y(_544__94_) );
INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_909_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf1), .B(clgen_enable_bF_buf7), .C(_707_), .Y(_910_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_910_), .Y(_911_) );
INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf0), .Y(_912_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_1702_), .C(_912__bF_buf5), .Y(_913_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_686__bF_buf8), .C(_913_), .Y(_914_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(wb_sel_i_3_bF_buf1_), .C(_711_), .Y(_915_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_915_), .C(_693__bF_buf3), .Y(_916_) );
OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(_693__bF_buf2), .C(_914_), .D(_916_), .Y(_544__93_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf0), .B(clgen_enable_bF_buf6), .C(_715_), .Y(_917_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_917_), .Y(_918_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_1867_), .C(_912__bF_buf3), .Y(_919_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_686__bF_buf7), .C(_919_), .Y(_920_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(wb_sel_i_3_bF_buf0_), .C(_719_), .Y(_921_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_921_), .C(_693__bF_buf1), .Y(_922_) );
OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_693__bF_buf0), .C(_920_), .D(_922_), .Y(_544__92_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf3), .B(clgen_enable_bF_buf5), .C(_722_), .Y(_923_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_923_), .Y(_924_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_1594_), .C(_912__bF_buf1), .Y(_925_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_686__bF_buf6), .C(_925_), .Y(_926_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(wb_sel_i_3_bF_buf6_), .C(_726_), .Y(_927_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_927_), .C(_693__bF_buf5), .Y(_928_) );
OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(_693__bF_buf4), .C(_926_), .D(_928_), .Y(_544__91_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf2), .B(clgen_enable_bF_buf4), .C(_729_), .Y(_929_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_929_), .Y(_930_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_1821_), .C(_912__bF_buf5), .Y(_931_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_686__bF_buf5), .C(_931_), .Y(_932_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(wb_sel_i_3_bF_buf5_), .C(_733_), .Y(_933_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_933_), .C(_693__bF_buf3), .Y(_934_) );
OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_693__bF_buf2), .C(_932_), .D(_934_), .Y(_544__90_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf1), .B(clgen_enable_bF_buf3), .C(_736_), .Y(_935_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_935_), .Y(_936_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_1688_), .C(_912__bF_buf3), .Y(_937_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_686__bF_buf4), .C(_937_), .Y(_938_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1688_), .B(wb_sel_i_3_bF_buf4_), .C(_740_), .Y(_939_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_939_), .C(_693__bF_buf1), .Y(_940_) );
OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1688_), .B(_693__bF_buf0), .C(_938_), .D(_940_), .Y(_544__89_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf0), .B(clgen_enable_bF_buf2), .C(_743_), .Y(_941_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_941_), .Y(_942_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_1912_), .C(_912__bF_buf1), .Y(_943_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_686__bF_buf3), .C(_943_), .Y(_944_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(wb_sel_i_3_bF_buf3_), .C(_747_), .Y(_945_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_945_), .C(_693__bF_buf5), .Y(_946_) );
OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_693__bF_buf4), .C(_944_), .D(_946_), .Y(_544__88_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf3), .B(clgen_enable_bF_buf1), .C(_751_), .Y(_947_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_909_), .Y(_948_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_948_), .C(_788__bF_buf4), .Y(_949_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_948_), .C(_949_), .Y(_950_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(wb_sel_i_2_bF_buf4_), .C(_755_), .Y(_951_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_951_), .C(_694__bF_buf7), .Y(_952_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_789__bF_buf1), .C(_950_), .D(_952_), .Y(_544__86_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf2), .B(clgen_enable_bF_buf0), .C(_758_), .Y(_953_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_953_), .Y(_954_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_1747_), .C(_912__bF_buf5), .Y(_955_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_686__bF_buf1), .C(_955_), .Y(_956_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(wb_sel_i_2_bF_buf3_), .C(_762_), .Y(_957_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_957_), .C(_693__bF_buf3), .Y(_958_) );
OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_693__bF_buf2), .C(_956_), .D(_958_), .Y(_544__85_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf1), .B(clgen_enable_bF_buf9), .C(_765_), .Y(_959_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_959_), .Y(_960_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_960_), .Y(_961_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .B(_961_), .C(_788__bF_buf3), .Y(_962_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_961_), .C(_962_), .Y(_963_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .B(wb_sel_i_2_bF_buf2_), .C(_769_), .Y(_964_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf0), .B(_964_), .C(_694__bF_buf6), .Y(_965_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .B(_789__bF_buf3), .C(_963_), .D(_965_), .Y(_544__84_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf0), .B(clgen_enable_bF_buf8), .C(_772_), .Y(_966_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_909_), .Y(_967_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1611_), .C(_912__bF_buf3), .Y(_968_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_686__bF_buf8), .C(_968_), .Y(_969_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(wb_sel_i_2_bF_buf1_), .C(_776_), .Y(_970_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_970_), .C(_693__bF_buf1), .Y(_971_) );
OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_693__bF_buf0), .C(_969_), .D(_971_), .Y(_544__83_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf3), .B(clgen_enable_bF_buf7), .C(_782_), .Y(_972_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_972_), .Y(_973_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_973_), .C(_788__bF_buf2), .Y(_974_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf7), .B(_973_), .C(_974_), .Y(_975_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(wb_sel_i_2_bF_buf0_), .C(_779_), .Y(_976_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_976_), .C(_694__bF_buf5), .Y(_977_) );
AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_789__bF_buf1), .C(_975_), .D(_977_), .Y(_544__82_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf2), .B(clgen_enable_bF_buf6), .C(_791_), .Y(_978_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_978_), .Y(_979_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_979_), .Y(_980_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_980_), .C(_788__bF_buf1), .Y(_981_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_980_), .C(_981_), .Y(_982_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(wb_sel_i_2_bF_buf6_), .C(_795_), .Y(_983_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf0), .B(_983_), .C(_694__bF_buf4), .Y(_984_) );
AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_789__bF_buf3), .C(_982_), .D(_984_), .Y(_544__81_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf1), .B(clgen_enable_bF_buf5), .C(_798_), .Y(_985_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_985_), .Y(_986_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_986_), .Y(_987_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_987_), .C(_788__bF_buf0), .Y(_988_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_987_), .C(_988_), .Y(_989_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(wb_sel_i_2_bF_buf5_), .C(_802_), .Y(_990_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_990_), .C(_694__bF_buf3), .Y(_991_) );
AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_789__bF_buf1), .C(_989_), .D(_991_), .Y(_544__80_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_2091__bF_buf3), .Y(_992_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_2025__bF_buf4), .B(_992_), .Y(_993_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_903_), .Y(_994_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_994_), .C(_788__bF_buf4), .Y(_995_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_994_), .C(_995_), .Y(_996_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(wb_sel_i_1_bF_buf3_), .C(_805_), .Y(_997_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf0), .B(_997_), .C(_694__bF_buf2), .Y(_998_) );
AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_789__bF_buf3), .C(_996_), .D(_998_), .Y(_544__78_) );
INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(_993_), .Y(_999_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_910_), .Y(_1000_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_1701_), .C(_912__bF_buf1), .Y(_1001_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_686__bF_buf3), .C(_1001_), .Y(_1002_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(wb_sel_i_1_bF_buf2_), .C(_821_), .Y(_1003_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1003_), .C(_693__bF_buf5), .Y(_1004_) );
OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_693__bF_buf4), .C(_1002_), .D(_1004_), .Y(_544__77_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_917_), .Y(_1005_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_1866_), .C(_912__bF_buf5), .Y(_1006_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_686__bF_buf2), .C(_1006_), .Y(_1007_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(wb_sel_i_1_bF_buf1_), .C(_827_), .Y(_1008_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_1008_), .C(_693__bF_buf3), .Y(_1009_) );
OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_693__bF_buf2), .C(_1007_), .D(_1009_), .Y(_544__76_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_923_), .Y(_1010_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1593_), .C(_912__bF_buf3), .Y(_1011_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_686__bF_buf1), .C(_1011_), .Y(_1012_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(wb_sel_i_1_bF_buf0_), .C(_833_), .Y(_1013_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_1013_), .C(_693__bF_buf1), .Y(_1014_) );
OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_693__bF_buf0), .C(_1012_), .D(_1014_), .Y(_544__75_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_929_), .Y(_1015_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1832_), .C(_912__bF_buf1), .Y(_1016_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_686__bF_buf0), .C(_1016_), .Y(_1017_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .B(wb_sel_i_1_bF_buf7_), .C(_836_), .Y(_1018_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1018_), .C(_693__bF_buf5), .Y(_1019_) );
OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .B(_693__bF_buf4), .C(_1017_), .D(_1019_), .Y(_544__74_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_935_), .Y(_1020_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1687_), .C(_912__bF_buf5), .Y(_1021_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_686__bF_buf8), .C(_1021_), .Y(_1022_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(wb_sel_i_1_bF_buf6_), .C(_849_), .Y(_1023_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_1023_), .C(_693__bF_buf3), .Y(_1024_) );
OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_693__bF_buf2), .C(_1022_), .D(_1024_), .Y(_544__73_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_941_), .Y(_1025_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1923_), .C(_912__bF_buf3), .Y(_1026_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_686__bF_buf7), .C(_1026_), .Y(_1027_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(wb_sel_i_1_bF_buf5_), .C(_855_), .Y(_1028_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_1028_), .C(_693__bF_buf1), .Y(_1029_) );
OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_693__bF_buf0), .C(_1027_), .D(_1029_), .Y(_544__72_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_947_), .Y(_1030_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1808_), .C(_912__bF_buf1), .Y(_1031_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_686__bF_buf6), .C(_1031_), .Y(_1032_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(wb_sel_i_0_bF_buf1_), .C(_861_), .Y(_1033_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1033_), .C(_693__bF_buf5), .Y(_1034_) );
OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(_693__bF_buf4), .C(_1032_), .D(_1034_), .Y(_544__70_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_953_), .Y(_1035_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1758_), .C(_912__bF_buf5), .Y(_1036_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_686__bF_buf5), .C(_1036_), .Y(_1037_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(wb_sel_i_0_bF_buf0_), .C(_867_), .Y(_1038_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_1038_), .C(_693__bF_buf3), .Y(_1039_) );
OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_693__bF_buf2), .C(_1037_), .D(_1039_), .Y(_544__69_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_960_), .Y(_1040_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(_1040_), .C(_788__bF_buf3), .Y(_1041_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1040_), .C(_1041_), .Y(_1042_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(wb_sel_i_0_bF_buf7_), .C(_873_), .Y(_1043_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_1043_), .C(_694__bF_buf1), .Y(_1044_) );
AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(_789__bF_buf1), .C(_1042_), .D(_1044_), .Y(_544__68_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_999_), .Y(_1045_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1618_), .C(_912__bF_buf3), .Y(_1046_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_686__bF_buf3), .C(_1046_), .Y(_1047_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(wb_sel_i_0_bF_buf6_), .C(_879_), .Y(_1048_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_1048_), .C(_693__bF_buf1), .Y(_1049_) );
OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_693__bF_buf0), .C(_1047_), .D(_1049_), .Y(_544__67_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_999_), .Y(_1050_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1855_), .C(_912__bF_buf1), .Y(_1051_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_686__bF_buf2), .C(_1051_), .Y(_1052_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(wb_sel_i_0_bF_buf5_), .C(_885_), .Y(_1053_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1053_), .C(_693__bF_buf5), .Y(_1054_) );
OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_693__bF_buf4), .C(_1052_), .D(_1054_), .Y(_544__66_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_999_), .Y(_1055_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1735_), .C(_912__bF_buf5), .Y(_1056_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_686__bF_buf1), .C(_1056_), .Y(_1057_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(wb_sel_i_0_bF_buf4_), .C(_891_), .Y(_1058_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_1058_), .C(_693__bF_buf3), .Y(_1059_) );
OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_693__bF_buf2), .C(_1057_), .D(_1059_), .Y(_544__65_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_986_), .Y(_1060_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1060_), .C(_788__bF_buf2), .Y(_1061_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_1060_), .C(_1061_), .Y(_1062_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(wb_sel_i_0_bF_buf3_), .C(_897_), .Y(_1063_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf0), .B(_1063_), .C(_694__bF_buf0), .Y(_1064_) );
AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_789__bF_buf3), .C(_1062_), .D(_1064_), .Y(_544__64_) );
INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(shift_latch_0_), .Y(_1065_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf4), .B(_1065_), .Y(_1066_) );
INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf6), .Y(_1067_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf7), .B(_2042_), .Y(_1068_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf1), .B(_902_), .Y(_1069_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1068_), .Y(_1070_) );
INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(shift_latch_1_), .Y(_1071_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf3), .B(_1071_), .Y(_1072_) );
INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf4), .Y(_1073_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1769_), .C(_1073__bF_buf4), .Y(_1074_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_686__bF_buf8), .C(_1074_), .Y(_1075_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(wb_sel_i_3_bF_buf2_), .C(_703_), .Y(_1076_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf3), .B(_1076_), .C(_1067__bF_buf6), .Y(_1077_) );
OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(_1067__bF_buf5), .C(_1075_), .D(_1077_), .Y(_544__62_) );
INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1078_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf0), .B(_910_), .Y(_1079_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1080_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1080_), .Y(_1081_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1707_), .C(_1073__bF_buf2), .Y(_1082_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_686__bF_buf7), .C(_1082_), .Y(_1083_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(wb_sel_i_3_bF_buf1_), .C(_711_), .Y(_1084_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf1), .B(_1084_), .C(_1067__bF_buf4), .Y(_1085_) );
OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_1067__bF_buf3), .C(_1083_), .D(_1085_), .Y(_544__61_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf4), .B(_917_), .Y(_1086_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_1086_), .Y(_1087_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1087_), .Y(_1088_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_1872_), .C(_1073__bF_buf0), .Y(_1089_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_686__bF_buf6), .C(_1089_), .Y(_1090_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(wb_sel_i_3_bF_buf0_), .C(_719_), .Y(_1091_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf4), .B(_1091_), .C(_1067__bF_buf2), .Y(_1092_) );
OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_1067__bF_buf1), .C(_1090_), .D(_1092_), .Y(_544__60_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf3), .B(_923_), .Y(_1093_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .Y(_1094_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1094_), .Y(_1095_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1571_), .C(_1073__bF_buf3), .Y(_1096_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_686__bF_buf5), .C(_1096_), .Y(_1097_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(wb_sel_i_3_bF_buf6_), .C(_726_), .Y(_1098_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf2), .B(_1098_), .C(_1067__bF_buf0), .Y(_1099_) );
OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1067__bF_buf6), .C(_1097_), .D(_1099_), .Y(_544__59_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf2), .B(_929_), .Y(_1100_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1100_), .Y(_1101_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1101_), .C(_1072__bF_buf3), .Y(_1102_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1101_), .C(_1102_), .Y(_1103_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(wb_sel_i_3_bF_buf5_), .C(_733_), .Y(_1104_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf2), .B(_1104_), .C(_1066__bF_buf5), .Y(_1105_) );
AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1066__bF_buf4), .C(_1103_), .D(_1105_), .Y(_544__58_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf1), .B(_935_), .Y(_1106_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_1106_), .Y(_1107_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1107_), .Y(_1108_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1683_), .C(_1073__bF_buf1), .Y(_1109_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_686__bF_buf3), .C(_1109_), .Y(_1110_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_1683_), .B(wb_sel_i_3_bF_buf4_), .C(_740_), .Y(_1111_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf0), .B(_1111_), .C(_1067__bF_buf5), .Y(_1112_) );
OAI22X1 OAI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1683_), .B(_1067__bF_buf4), .C(_1110_), .D(_1112_), .Y(_544__57_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf0), .B(_941_), .Y(_1113_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .Y(_1114_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1114_), .Y(_1115_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1907_), .C(_1073__bF_buf4), .Y(_1116_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_686__bF_buf2), .C(_1116_), .Y(_1117_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(wb_sel_i_3_bF_buf3_), .C(_747_), .Y(_1118_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf3), .B(_1118_), .C(_1067__bF_buf3), .Y(_1119_) );
OAI22X1 OAI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_1067__bF_buf2), .C(_1117_), .D(_1119_), .Y(_544__56_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf4), .B(_947_), .Y(_1120_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_1068_), .Y(_1121_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1792_), .C(_1073__bF_buf2), .Y(_1122_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_686__bF_buf1), .C(_1122_), .Y(_1123_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(wb_sel_i_2_bF_buf4_), .C(_755_), .Y(_1124_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf1), .B(_1124_), .C(_1067__bF_buf1), .Y(_1125_) );
OAI22X1 OAI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1067__bF_buf0), .C(_1123_), .D(_1125_), .Y(_544__54_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf3), .B(_953_), .Y(_1126_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1126_), .B(_1068_), .Y(_1127_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1742_), .C(_1073__bF_buf0), .Y(_1128_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_686__bF_buf0), .C(_1128_), .Y(_1129_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(wb_sel_i_2_bF_buf3_), .C(_762_), .Y(_1130_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf4), .B(_1130_), .C(_1067__bF_buf6), .Y(_1131_) );
OAI22X1 OAI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(_1067__bF_buf5), .C(_1129_), .D(_1131_), .Y(_544__53_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf2), .B(_691_), .C(_960_), .Y(_1132_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .Y(_1133_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1133_), .Y(_1134_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1134_), .C(_1072__bF_buf1), .Y(_1135_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_1134_), .C(_1135_), .Y(_1136_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(wb_sel_i_2_bF_buf2_), .C(_769_), .Y(_1137_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf0), .B(_1137_), .C(_1066__bF_buf3), .Y(_1138_) );
AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1066__bF_buf2), .C(_1136_), .D(_1138_), .Y(_544__52_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf2), .B(_966_), .Y(_1139_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1068_), .Y(_1140_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1605_), .C(_1073__bF_buf3), .Y(_1141_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_686__bF_buf7), .C(_1141_), .Y(_1142_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .B(wb_sel_i_2_bF_buf1_), .C(_776_), .Y(_1143_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf2), .B(_1143_), .C(_1067__bF_buf4), .Y(_1144_) );
OAI22X1 OAI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .B(_1067__bF_buf3), .C(_1142_), .D(_1144_), .Y(_544__51_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf1), .B(_972_), .Y(_1145_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1145_), .Y(_1146_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1146_), .C(_1072__bF_buf4), .Y(_1147_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_1146_), .C(_1147_), .Y(_1148_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(wb_sel_i_2_bF_buf0_), .C(_779_), .Y(_1149_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf3), .B(_1149_), .C(_1066__bF_buf1), .Y(_1150_) );
AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1066__bF_buf0), .C(_1148_), .D(_1150_), .Y(_544__50_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf1), .B(_691_), .C(_979_), .Y(_1151_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1151_), .Y(_1152_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_1724_), .C(_1073__bF_buf1), .Y(_1153_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_686__bF_buf5), .C(_1153_), .Y(_1154_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(wb_sel_i_2_bF_buf6_), .C(_795_), .Y(_1155_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf0), .B(_1155_), .C(_1067__bF_buf2), .Y(_1156_) );
OAI22X1 OAI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_1067__bF_buf1), .C(_1154_), .D(_1156_), .Y(_544__49_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf0), .B(_985_), .Y(_1157_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1157_), .Y(_1158_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1158_), .C(_1072__bF_buf2), .Y(_1159_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1158_), .C(_1159_), .Y(_1160_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(wb_sel_i_2_bF_buf5_), .C(_802_), .Y(_1161_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf1), .B(_1161_), .C(_1066__bF_buf6), .Y(_1162_) );
AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1066__bF_buf5), .C(_1160_), .D(_1162_), .Y(_544__48_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf6), .B(_808_), .Y(_1163_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1069_), .Y(_1164_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1164_), .C(_1072__bF_buf0), .Y(_1165_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_1164_), .C(_1165_), .Y(_1166_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(wb_sel_i_1_bF_buf4_), .C(_805_), .Y(_1167_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf4), .B(_1167_), .C(_1066__bF_buf4), .Y(_1168_) );
AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1066__bF_buf3), .C(_1166_), .D(_1168_), .Y(_544__46_) );
INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .Y(_1169_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1080_), .Y(_1170_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1706_), .C(_1073__bF_buf4), .Y(_1171_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_686__bF_buf2), .C(_1171_), .Y(_1172_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(wb_sel_i_1_bF_buf3_), .C(_821_), .Y(_1173_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf3), .B(_1173_), .C(_1067__bF_buf0), .Y(_1174_) );
OAI22X1 OAI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1067__bF_buf6), .C(_1172_), .D(_1174_), .Y(_544__45_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1087_), .Y(_1175_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1871_), .C(_1073__bF_buf2), .Y(_1176_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_686__bF_buf1), .C(_1176_), .Y(_1177_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_1871_), .B(wb_sel_i_1_bF_buf2_), .C(_827_), .Y(_1178_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf1), .B(_1178_), .C(_1067__bF_buf5), .Y(_1179_) );
OAI22X1 OAI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1871_), .B(_1067__bF_buf4), .C(_1177_), .D(_1179_), .Y(_544__44_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1094_), .Y(_1180_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_1570_), .C(_1073__bF_buf0), .Y(_1181_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_686__bF_buf0), .C(_1181_), .Y(_1182_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(wb_sel_i_1_bF_buf1_), .C(_833_), .Y(_1183_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf4), .B(_1183_), .C(_1067__bF_buf3), .Y(_1184_) );
OAI22X1 OAI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1067__bF_buf2), .C(_1182_), .D(_1184_), .Y(_544__43_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1100_), .Y(_1185_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1185_), .C(_1072__bF_buf3), .Y(_1186_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_1185_), .C(_1186_), .Y(_1187_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(wb_sel_i_1_bF_buf0_), .C(_836_), .Y(_1188_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf2), .B(_1188_), .C(_1066__bF_buf2), .Y(_1189_) );
AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1066__bF_buf1), .C(_1187_), .D(_1189_), .Y(_544__42_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1107_), .Y(_1190_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1682_), .C(_1073__bF_buf3), .Y(_1191_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_686__bF_buf7), .C(_1191_), .Y(_1192_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(wb_sel_i_1_bF_buf7_), .C(_849_), .Y(_1193_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf2), .B(_1193_), .C(_1067__bF_buf1), .Y(_1194_) );
OAI22X1 OAI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(_1067__bF_buf0), .C(_1192_), .D(_1194_), .Y(_544__41_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1114_), .Y(_1195_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1918_), .C(_1073__bF_buf1), .Y(_1196_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_686__bF_buf6), .C(_1196_), .Y(_1197_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(wb_sel_i_1_bF_buf6_), .C(_855_), .Y(_1198_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf0), .B(_1198_), .C(_1067__bF_buf6), .Y(_1199_) );
OAI22X1 OAI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(_1067__bF_buf5), .C(_1197_), .D(_1199_), .Y(_544__40_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1120_), .Y(_1200_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1200_), .C(_1072__bF_buf1), .Y(_1201_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_1200_), .C(_1201_), .Y(_1202_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(wb_sel_i_0_bF_buf2_), .C(_861_), .Y(_1203_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf0), .B(_1203_), .C(_1066__bF_buf0), .Y(_1204_) );
AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1066__bF_buf6), .C(_1202_), .D(_1204_), .Y(_544__38_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1126_), .Y(_1205_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1205_), .C(_1072__bF_buf4), .Y(_1206_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1205_), .C(_1206_), .Y(_1207_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(wb_sel_i_0_bF_buf1_), .C(_867_), .Y(_1208_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf3), .B(_1208_), .C(_1066__bF_buf5), .Y(_1209_) );
AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1066__bF_buf4), .C(_1207_), .D(_1209_), .Y(_544__37_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1133_), .Y(_1210_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(_1210_), .C(_1072__bF_buf2), .Y(_1211_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_1210_), .C(_1211_), .Y(_1212_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(wb_sel_i_0_bF_buf0_), .C(_873_), .Y(_1213_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf1), .B(_1213_), .C(_1066__bF_buf3), .Y(_1214_) );
AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(_1066__bF_buf2), .C(_1212_), .D(_1214_), .Y(_544__36_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1139_), .Y(_1215_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1215_), .C(_1072__bF_buf0), .Y(_1216_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_1215_), .C(_1216_), .Y(_1217_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(wb_sel_i_0_bF_buf7_), .C(_879_), .Y(_1218_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf4), .B(_1218_), .C(_1066__bF_buf1), .Y(_1219_) );
AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1066__bF_buf0), .C(_1217_), .D(_1219_), .Y(_544__35_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1145_), .Y(_1220_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1220_), .C(_1072__bF_buf3), .Y(_1221_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf1), .B(_1220_), .C(_1221_), .Y(_1222_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(wb_sel_i_0_bF_buf6_), .C(_885_), .Y(_1223_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf2), .B(_1223_), .C(_1066__bF_buf6), .Y(_1224_) );
AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1066__bF_buf5), .C(_1222_), .D(_1224_), .Y(_544__34_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1151_), .Y(_1225_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1730_), .C(_1073__bF_buf4), .Y(_1226_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_686__bF_buf0), .C(_1226_), .Y(_1227_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(wb_sel_i_0_bF_buf5_), .C(_891_), .Y(_1228_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_1073__bF_buf3), .B(_1228_), .C(_1067__bF_buf4), .Y(_1229_) );
OAI22X1 OAI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1067__bF_buf3), .C(_1227_), .D(_1229_), .Y(_544__33_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1157_), .Y(_1230_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1230_), .C(_1072__bF_buf1), .Y(_1231_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf8), .B(_1230_), .C(_1231_), .Y(_1232_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(wb_sel_i_0_bF_buf4_), .C(_897_), .Y(_1233_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf0), .B(_1233_), .C(_1066__bF_buf4), .Y(_1234_) );
AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1066__bF_buf3), .C(_1232_), .D(_1234_), .Y(_544__32_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[30]), .B(rx_30_), .S(wb_sel_i_3_bF_buf2_), .Y(_1235_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf5), .B(_900_), .Y(_1236_) );
INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .Y(_1237_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf0), .B(_1071_), .C(_1069_), .Y(_1238_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1238_), .Y(_1239_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf0), .B(_1772_), .S(_1239_), .Y(_1240_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_1065_), .C(_1240_), .Y(_1241_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1235_), .C(_1241_), .Y(_544__30_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[29]), .B(rx_29_), .S(wb_sel_i_3_bF_buf1_), .Y(_1242_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf8), .B(_1071_), .C(_1079_), .Y(_1243_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1243_), .Y(_1244_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1711_), .S(_1244_), .Y(_1245_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf7), .B(_1065_), .C(_1245_), .Y(_1246_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1242_), .C(_1246_), .Y(_544__29_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[28]), .B(rx_28_), .S(wb_sel_i_3_bF_buf0_), .Y(_1247_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf6), .B(_1071_), .C(_1086_), .Y(_1248_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1248_), .Y(_1249_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf3), .B(_1876_), .S(_1249_), .Y(_1250_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf5), .B(_1065_), .C(_1250_), .Y(_1251_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf0), .B(_1247_), .C(_1251_), .Y(_544__28_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_1584_), .B(wb_sel_i_3_bF_buf6_), .C(_726_), .Y(_1252_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf2), .B(_1252_), .Y(_1253_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf4), .B(_1071_), .C(_1093_), .Y(_1254_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1254_), .Y(_1255_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf2), .B(_1255_), .Y(_1256_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(rx_27_), .C(_1067__bF_buf6), .Y(_1257_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1257_), .C(_1253_), .Y(_544__27_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[26]), .B(rx_26_), .S(wb_sel_i_3_bF_buf5_), .Y(_1258_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf3), .B(_1071_), .C(_1100_), .Y(_1259_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1259_), .Y(_1260_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1819_), .S(_1260_), .Y(_1261_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf2), .B(_1065_), .C(_1261_), .Y(_1262_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1258_), .C(_1262_), .Y(_544__26_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf1), .B(_1071_), .C(_1106_), .Y(_1263_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1263_), .Y(_1264_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_685__bF_buf0), .Y(_1265_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(rx_25_), .B(_1264_), .C(_1265_), .Y(_1266_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[25]), .B(rx_25_), .S(wb_sel_i_3_bF_buf4_), .Y(_1267_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1267_), .S(_1067__bF_buf4), .Y(_544__25_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[24]), .B(rx_24_), .S(wb_sel_i_3_bF_buf3_), .Y(_1268_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf0), .B(_1071_), .C(_1113_), .Y(_1269_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1269_), .Y(_1270_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1910_), .S(_1270_), .Y(_1271_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_1065_), .C(_1271_), .Y(_1272_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1268_), .C(_1272_), .Y(_544__24_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[22]), .B(rx_22_), .S(wb_sel_i_2_bF_buf4_), .Y(_1273_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf8), .B(_1071_), .C(_1120_), .Y(_1274_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1274_), .Y(_1275_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf3), .B(_1795_), .S(_1275_), .Y(_1276_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf7), .B(_1065_), .C(_1276_), .Y(_1277_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1273_), .C(_1277_), .Y(_544__22_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(wb_sel_i_2_bF_buf3_), .C(_762_), .Y(_1278_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf1), .B(_1278_), .Y(_1279_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf6), .B(_1071_), .C(_1126_), .Y(_1280_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1280_), .Y(_1281_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf2), .B(_1281_), .Y(_1282_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_1281_), .B(rx_21_), .C(_1067__bF_buf1), .Y(_1283_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1283_), .C(_1279_), .Y(_544__21_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(wb_sel_i_2_bF_buf2_), .C(_769_), .Y(_1284_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf0), .B(_1284_), .Y(_1285_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf5), .B(_1071_), .C(_1133_), .Y(_1286_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1286_), .Y(_1287_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1287_), .Y(_1288_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(rx_20_), .C(_1067__bF_buf0), .Y(_1289_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_1288_), .B(_1289_), .C(_1285_), .Y(_544__20_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(wb_sel_i_2_bF_buf1_), .C(_776_), .Y(_1290_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf6), .B(_1290_), .Y(_1291_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf4), .B(_1071_), .C(_1139_), .Y(_1292_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1292_), .Y(_1293_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_685__bF_buf0), .Y(_1294_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(rx_19_), .B(_1293_), .C(_1294_), .Y(_1295_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1066__bF_buf5), .C(_1291_), .Y(_544__19_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(wb_sel_i_2_bF_buf0_), .C(_779_), .Y(_1296_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf4), .B(_1296_), .Y(_1297_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf3), .B(_1071_), .C(_1145_), .Y(_1298_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1298_), .Y(_1299_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1299_), .Y(_1300_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(rx_18_), .C(_1067__bF_buf6), .Y(_1301_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1301_), .C(_1297_), .Y(_544__18_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(wb_sel_i_2_bF_buf6_), .C(_795_), .Y(_1302_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf3), .B(_1302_), .Y(_1303_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf4), .B(_1151_), .Y(_1304_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1304_), .Y(_1305_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_686__bF_buf7), .Y(_1306_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .Y(_1307_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(rx_17_), .C(_1067__bF_buf5), .Y(_1308_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1308_), .C(_1303_), .Y(_544__17_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(wb_sel_i_2_bF_buf5_), .C(_802_), .Y(_1309_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf2), .B(_1309_), .Y(_1310_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf2), .B(_1071_), .C(_1157_), .Y(_1311_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1311_), .Y(_1312_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_685__bF_buf3), .Y(_1313_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(rx_16_), .B(_1312_), .C(_1313_), .Y(_1314_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1066__bF_buf1), .C(_1310_), .Y(_544__16_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[14]), .B(rx_14_), .S(wb_sel_i_1_bF_buf5_), .Y(_1315_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_2078__bF_buf4), .B(_992_), .Y(_1316_) );
INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .Y(_1317_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1238_), .Y(_1318_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf2), .B(_1783_), .S(_1318_), .Y(_1319_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf1), .B(_1065_), .C(_1319_), .Y(_1320_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1315_), .C(_1320_), .Y(_544__14_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_1710_), .B(wb_sel_i_1_bF_buf4_), .C(_821_), .Y(_1321_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf0), .B(_1321_), .Y(_1322_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1243_), .Y(_1323_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1323_), .Y(_1324_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(rx_13_), .C(_1067__bF_buf3), .Y(_1325_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_1325_), .C(_1322_), .Y(_544__13_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[12]), .B(rx_12_), .S(wb_sel_i_1_bF_buf3_), .Y(_1326_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1248_), .Y(_1327_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf0), .B(_1875_), .S(_1327_), .Y(_1328_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf0), .B(_1065_), .C(_1328_), .Y(_1329_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1326_), .C(_1329_), .Y(_544__12_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .B(wb_sel_i_1_bF_buf2_), .C(_833_), .Y(_1330_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf6), .B(_1330_), .Y(_1331_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1254_), .Y(_1332_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1332_), .Y(_1333_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(rx_11_), .C(_1067__bF_buf1), .Y(_1334_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1334_), .C(_1331_), .Y(_544__11_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(wb_sel_i_1_bF_buf1_), .C(_836_), .Y(_1335_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf5), .B(_1335_), .Y(_1336_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1259_), .Y(_1337_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf3), .B(_1337_), .Y(_1338_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_1337_), .B(rx_10_), .C(_1067__bF_buf0), .Y(_1339_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1339_), .C(_1336_), .Y(_544__10_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .B(wb_sel_i_1_bF_buf0_), .C(_849_), .Y(_1340_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf4), .B(_1340_), .Y(_1341_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1263_), .Y(_1342_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf2), .B(_1342_), .Y(_1343_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(rx_9_), .C(_1067__bF_buf6), .Y(_1344_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1344_), .C(_1341_), .Y(_544__9_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(wb_sel_i_1_bF_buf7_), .C(_855_), .Y(_1345_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf3), .B(_1345_), .Y(_1346_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1269_), .Y(_1347_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1347_), .Y(_1348_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(rx_8_), .C(_1067__bF_buf5), .Y(_1349_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1349_), .C(_1346_), .Y(_544__8_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[6]), .B(rx_6_), .S(wb_sel_i_0_bF_buf3_), .Y(_1350_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1274_), .Y(_1351_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf0), .B(_1806_), .S(_1351_), .Y(_1352_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_1065_), .C(_1352_), .Y(_1353_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1350_), .C(_1353_), .Y(_544__6_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[5]), .B(rx_5_), .S(wb_sel_i_0_bF_buf2_), .Y(_1354_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1280_), .Y(_1355_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1756_), .S(_1355_), .Y(_1356_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf8), .B(_1065_), .C(_1356_), .Y(_1357_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf3), .B(_1354_), .C(_1357_), .Y(_544__5_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(wb_sel_i_0_bF_buf1_), .C(_873_), .Y(_1358_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf2), .B(_1358_), .Y(_1359_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1286_), .Y(_1360_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_685__bF_buf3), .Y(_1361_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(rx_4_), .B(_1360_), .C(_1361_), .Y(_1362_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1066__bF_buf1), .C(_1359_), .Y(_544__4_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[3]), .B(rx_3_), .S(wb_sel_i_0_bF_buf0_), .Y(_1363_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1292_), .Y(_1364_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf2), .B(_1616_), .S(_1364_), .Y(_1365_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf7), .B(_1065_), .C(_1365_), .Y(_1366_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf2), .B(_1363_), .C(_1366_), .Y(_544__3_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[2]), .B(rx_2_), .S(wb_sel_i_0_bF_buf7_), .Y(_1367_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1298_), .Y(_1368_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1853_), .S(_1368_), .Y(_1369_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf6), .B(_1065_), .C(_1369_), .Y(_1370_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf1), .B(_1367_), .C(_1370_), .Y(_544__2_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(wb_sel_i_0_bF_buf6_), .C(_891_), .Y(_1371_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf0), .B(_1371_), .Y(_1372_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1304_), .Y(_1373_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_686__bF_buf6), .Y(_1374_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .Y(_1375_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(rx_1_), .C(_1067__bF_buf0), .Y(_1376_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_1376_), .C(_1372_), .Y(_544__1_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[0]), .B(rx_0_), .S(wb_sel_i_0_bF_buf5_), .Y(_1377_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1311_), .Y(_1378_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf0), .B(_1944_), .S(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf5), .B(_1065_), .C(_1379_), .Y(_1380_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf6), .B(_1377_), .C(_1380_), .Y(_544__0_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf0), .B(clgen_enable_bF_buf4), .C(_2071_), .Y(_1381_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_1381_), .Y(_1382_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1632_), .C(_912__bF_buf3), .Y(_1383_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_686__bF_buf5), .C(_1383_), .Y(_1384_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(wb_sel_i_3_bF_buf2_), .C(_695_), .Y(_1385_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(_1385_), .C(_693__bF_buf1), .Y(_1386_) );
OAI22X1 OAI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_693__bF_buf0), .C(_1384_), .D(_1386_), .Y(_544__95_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_809_), .Y(_1387_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1387_), .C(_688__bF_buf5), .Y(_1388_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1387_), .C(_1388_), .Y(_1389_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_1_bF_buf6_), .B(wb_dat_i[15]), .Y(_1390_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(wb_sel_i_1_bF_buf5_), .C(_1390_), .Y(_1391_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf4), .B(_1391_), .C(_694__bF_buf7), .Y(_1392_) );
AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_694__bF_buf6), .C(_1389_), .D(_1392_), .Y(_544__111_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_750_), .Y(_1393_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_1393_), .Y(_1394_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1394_), .C(_688__bF_buf3), .Y(_1395_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf3), .B(_1394_), .C(_1395_), .Y(_1396_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_2_bF_buf4_), .B(wb_dat_i[23]), .Y(_1397_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(wb_sel_i_2_bF_buf3_), .C(_1397_), .Y(_1398_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf2), .B(_1398_), .C(_694__bF_buf5), .Y(_1399_) );
AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_694__bF_buf4), .C(_1396_), .D(_1399_), .Y(_544__119_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf4), .B(_1381_), .Y(_1400_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1400_), .Y(_1401_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1401_), .C(_1072__bF_buf3), .Y(_1402_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf2), .B(_1401_), .C(_1402_), .Y(_1403_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(wb_sel_i_3_bF_buf1_), .C(_695_), .Y(_1404_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf2), .B(_1404_), .C(_1066__bF_buf6), .Y(_1405_) );
AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1066__bF_buf5), .C(_1403_), .D(_1405_), .Y(_544__63_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1381_), .Y(_1406_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1643_), .C(_912__bF_buf1), .Y(_1407_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_686__bF_buf1), .C(_1407_), .Y(_1408_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(wb_sel_i_1_bF_buf4_), .C(_1390_), .Y(_1409_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1409_), .C(_693__bF_buf5), .Y(_1410_) );
OAI22X1 OAI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_693__bF_buf4), .C(_1408_), .D(_1410_), .Y(_544__79_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_687__bF_buf3), .B(clgen_enable_bF_buf3), .C(_1393_), .Y(_1411_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_909_), .Y(_1412_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1412_), .C(_788__bF_buf3), .Y(_1413_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf0), .B(_1412_), .C(_1413_), .Y(_1414_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(wb_sel_i_2_bF_buf2_), .C(_1397_), .Y(_1415_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_789__bF_buf2), .B(_1415_), .C(_694__bF_buf3), .Y(_1416_) );
AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_789__bF_buf1), .C(_1414_), .D(_1416_), .Y(_544__87_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1411_), .Y(_1417_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1671_), .C(_912__bF_buf5), .Y(_1418_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_686__bF_buf8), .C(_1418_), .Y(_1419_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(wb_sel_i_0_bF_buf4_), .B(wb_dat_i[7]), .Y(_1420_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(wb_sel_i_0_bF_buf3_), .C(_1420_), .Y(_1421_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_1421_), .C(_693__bF_buf3), .Y(_1422_) );
OAI22X1 OAI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_693__bF_buf2), .C(_1419_), .D(_1422_), .Y(_544__71_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[31]), .B(rx_31_), .S(wb_sel_i_3_bF_buf0_), .Y(_1423_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf2), .B(_1071_), .C(_1400_), .Y(_1424_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1424_), .Y(_1425_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf4), .B(_1630_), .S(_1425_), .Y(_1426_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf1), .B(_1065_), .C(_1426_), .Y(_1427_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf5), .B(_1423_), .C(_1427_), .Y(_544__31_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1400_), .Y(_1428_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1428_), .C(_1072__bF_buf1), .Y(_1429_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf7), .B(_1428_), .C(_1429_), .Y(_1430_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(wb_sel_i_1_bF_buf3_), .C(_1390_), .Y(_1431_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf0), .B(_1431_), .C(_1066__bF_buf4), .Y(_1432_) );
AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1066__bF_buf3), .C(_1430_), .D(_1432_), .Y(_544__47_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_788__bF_buf2), .B(_1411_), .Y(_1433_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1433_), .Y(_1434_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1434_), .C(_1072__bF_buf4), .Y(_1435_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf6), .B(_1434_), .C(_1435_), .Y(_1436_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(wb_sel_i_2_bF_buf1_), .C(_1397_), .Y(_1437_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf3), .B(_1437_), .C(_1066__bF_buf2), .Y(_1438_) );
AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1066__bF_buf1), .C(_1436_), .D(_1438_), .Y(_544__55_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1433_), .Y(_1439_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1439_), .C(_1072__bF_buf2), .Y(_1440_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf5), .B(_1439_), .C(_1440_), .Y(_1441_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(wb_sel_i_0_bF_buf2_), .C(_1420_), .Y(_1442_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1072__bF_buf1), .B(_1442_), .C(_1066__bF_buf0), .Y(_1443_) );
AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1066__bF_buf6), .C(_1441_), .D(_1443_), .Y(_544__39_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_1393_), .Y(_1444_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(_1444_), .C(_688__bF_buf1), .Y(_1445_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_686__bF_buf4), .B(_1444_), .C(_1445_), .Y(_1446_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(wb_sel_i_0_bF_buf1_), .C(_1420_), .Y(_1447_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_688__bF_buf0), .B(_1447_), .C(_694__bF_buf2), .Y(_1448_) );
AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(_694__bF_buf1), .C(_1446_), .D(_1448_), .Y(_544__103_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(wb_sel_i_1_bF_buf2_), .C(_1390_), .Y(_1449_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf5), .B(_1449_), .Y(_1450_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1424_), .Y(_1451_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_685__bF_buf3), .Y(_1452_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(rx_15_), .B(_1451_), .C(_1452_), .Y(_1453_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1066__bF_buf4), .C(_1450_), .Y(_544__15_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_1658_), .B(wb_sel_i_2_bF_buf0_), .C(_1397_), .Y(_1454_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1066__bF_buf3), .B(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf0), .B(_1071_), .C(_1433_), .Y(_1456_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1456_), .Y(_1457_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .B(_685__bF_buf2), .Y(_1458_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(rx_23_), .B(_1457_), .C(_1458_), .Y(_1459_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1066__bF_buf2), .C(_1455_), .Y(_544__23_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(wb_dat_i[7]), .B(rx_7_), .S(wb_sel_i_0_bF_buf0_), .Y(_1460_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1456_), .Y(_1461_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_685__bF_buf1), .B(_1669_), .S(_1461_), .Y(_1462_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(_1065_), .C(_1462_), .Y(_1463_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_1067__bF_buf4), .B(_1460_), .C(_1463_), .Y(_544__7_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_0_), .B(clgen_pos_edge), .Y(_1464_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .B(clgen_enable_bF_buf8), .Y(_1465_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf7), .B(_1464_), .C(_1465_), .Y(_543__0_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_1510_), .Y(_1466_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_1_), .B(clgen_pos_edge), .C(clgen_enable_bF_buf6), .Y(_1467_) );
OAI22X1 OAI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(clgen_enable_bF_buf5), .C(_1466_), .D(_1467_), .Y(_543__1_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_1519_), .Y(_1468_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_2_), .B(clgen_pos_edge), .C(clgen_enable_bF_buf4), .Y(_1469_) );
OAI22X1 OAI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(clgen_enable_bF_buf3), .C(_1468_), .D(_1469_), .Y(_543__2_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(clgen_pos_edge), .B(_1535_), .Y(_1470_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_3_), .B(clgen_pos_edge), .C(_1470_), .Y(_1471_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(char_len_3_), .B(_692_), .Y(_1472_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_692_), .C(_1472_), .Y(_543__3_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(clgen_pos_edge), .B(_1574_), .Y(_1473_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_4_), .B(clgen_pos_edge), .C(_1473_), .Y(_1474_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .B(_692_), .Y(_1475_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_692_), .C(_1475_), .Y(_543__4_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_1567_), .Y(_1476_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_5_), .B(clgen_pos_edge), .C(clgen_enable_bF_buf2), .Y(_1477_) );
OAI22X1 OAI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(clgen_enable_bF_buf1), .C(_1476_), .D(_1477_), .Y(_543__5_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(char_len_6_), .Y(_1478_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_2140_), .C(shift_cnt_6_), .Y(_1479_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_1498_), .Y(_1480_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_1480_), .Y(_1481_) );
AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_692_), .C(_1481_), .D(_1479_), .Y(_543__6_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_7_), .B(clgen_enable_bF_buf0), .Y(_1482_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .B(char_len_4_), .Y(_1483_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1551_), .C(_1483_), .Y(_1484_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1521_), .C(_1465_), .Y(_1485_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_1484_), .Y(_1486_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(shift_cnt_7_), .B(_692_), .Y(_1487_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_1480_), .C(_1486_), .Y(_1488_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1482_), .C(_1488_), .Y(_543__7_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(clgen_enable_bF_buf9), .B(clgen_go), .Y(_1489_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_1480_), .C(_1489_), .Y(_546_) );
INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(wb_rst_i), .Y(_547_) );
DFFSR DFFSR_116 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf0), .D(_544__0_), .Q(rx_0_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_117 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf0), .D(_544__1_), .Q(rx_1_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_118 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf0), .D(_544__2_), .Q(rx_2_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_119 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__3_), .Q(rx_3_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_120 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__4_), .Q(rx_4_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_121 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf3), .D(_544__5_), .Q(rx_5_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_122 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf3), .D(_544__6_), .Q(rx_6_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_123 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf3), .D(_544__7_), .Q(rx_7_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_124 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf3), .D(_544__8_), .Q(rx_8_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_125 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf3), .D(_544__9_), .Q(rx_9_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_126 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf3), .D(_544__10_), .Q(rx_10_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_127 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf3), .D(_544__11_), .Q(rx_11_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_128 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf3), .D(_544__12_), .Q(rx_12_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_129 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf3), .D(_544__13_), .Q(rx_13_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_130 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf3), .D(_544__14_), .Q(rx_14_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_131 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf3), .D(_544__15_), .Q(rx_15_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_132 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf3), .D(_544__16_), .Q(rx_16_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_133 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf3), .D(_544__17_), .Q(rx_17_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_134 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__18_), .Q(rx_18_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_135 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__19_), .Q(rx_19_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_136 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf2), .D(_544__20_), .Q(rx_20_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_137 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf2), .D(_544__21_), .Q(rx_21_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_138 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf2), .D(_544__22_), .Q(rx_22_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_139 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf2), .D(_544__23_), .Q(rx_23_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_140 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf2), .D(_544__24_), .Q(rx_24_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_141 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf2), .D(_544__25_), .Q(rx_25_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_142 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf2), .D(_544__26_), .Q(rx_26_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_143 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf2), .D(_544__27_), .Q(rx_27_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_144 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf2), .D(_544__28_), .Q(rx_28_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_145 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf2), .D(_544__29_), .Q(rx_29_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_146 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf2), .D(_544__30_), .Q(rx_30_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_147 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf2), .D(_544__31_), .Q(rx_31_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_148 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf2), .D(_544__32_), .Q(rx_32_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_149 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__33_), .Q(rx_33_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_150 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__34_), .Q(rx_34_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_151 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf1), .D(_544__35_), .Q(rx_35_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_152 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf1), .D(_544__36_), .Q(rx_36_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_153 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf1), .D(_544__37_), .Q(rx_37_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_154 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf1), .D(_544__38_), .Q(rx_38_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_155 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf1), .D(_544__39_), .Q(rx_39_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_156 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf1), .D(_544__40_), .Q(rx_40_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_157 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf1), .D(_544__41_), .Q(rx_41_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_158 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf1), .D(_544__42_), .Q(rx_42_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_159 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf1), .D(_544__43_), .Q(rx_43_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_160 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf1), .D(_544__44_), .Q(rx_44_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_161 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf1), .D(_544__45_), .Q(rx_45_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_162 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf1), .D(_544__46_), .Q(rx_46_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_163 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf1), .D(_544__47_), .Q(rx_47_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_164 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__48_), .Q(rx_48_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_165 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__49_), .Q(rx_49_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_166 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf0), .D(_544__50_), .Q(rx_50_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_167 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf0), .D(_544__51_), .Q(rx_51_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_168 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf0), .D(_544__52_), .Q(rx_52_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_169 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf0), .D(_544__53_), .Q(rx_53_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_170 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf0), .D(_544__54_), .Q(rx_54_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_171 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf0), .D(_544__55_), .Q(rx_55_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_172 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf0), .D(_544__56_), .Q(rx_56_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_173 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf0), .D(_544__57_), .Q(rx_57_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_174 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf0), .D(_544__58_), .Q(rx_58_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_175 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf0), .D(_544__59_), .Q(rx_59_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_176 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf0), .D(_544__60_), .Q(rx_60_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_177 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf0), .D(_544__61_), .Q(rx_61_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_178 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf0), .D(_544__62_), .Q(rx_62_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_179 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__63_), .Q(rx_63_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_180 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__64_), .Q(rx_64_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_181 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf3), .D(_544__65_), .Q(rx_65_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_182 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf3), .D(_544__66_), .Q(rx_66_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_183 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf3), .D(_544__67_), .Q(rx_67_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_184 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf3), .D(_544__68_), .Q(rx_68_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_185 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf3), .D(_544__69_), .Q(rx_69_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_186 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf3), .D(_544__70_), .Q(rx_70_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_187 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf3), .D(_544__71_), .Q(rx_71_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_188 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf3), .D(_544__72_), .Q(rx_72_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_189 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf3), .D(_544__73_), .Q(rx_73_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_190 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf3), .D(_544__74_), .Q(rx_74_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_191 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf3), .D(_544__75_), .Q(rx_75_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_192 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf3), .D(_544__76_), .Q(rx_76_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_193 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf3), .D(_544__77_), .Q(rx_77_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_194 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__78_), .Q(rx_78_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_195 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__79_), .Q(rx_79_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_196 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf2), .D(_544__80_), .Q(rx_80_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_197 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf2), .D(_544__81_), .Q(rx_81_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_198 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf2), .D(_544__82_), .Q(rx_82_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_199 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf2), .D(_544__83_), .Q(rx_83_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_200 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf2), .D(_544__84_), .Q(rx_84_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_201 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf2), .D(_544__85_), .Q(rx_85_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_202 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf2), .D(_544__86_), .Q(rx_86_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_203 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf2), .D(_544__87_), .Q(rx_87_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_204 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf2), .D(_544__88_), .Q(rx_88_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_205 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf2), .D(_544__89_), .Q(rx_89_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_206 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf2), .D(_544__90_), .Q(rx_90_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_207 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf2), .D(_544__91_), .Q(rx_91_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_208 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf2), .D(_544__92_), .Q(rx_92_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_209 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__93_), .Q(rx_93_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_210 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__94_), .Q(rx_94_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_211 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf1), .D(_544__95_), .Q(rx_95_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_212 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf1), .D(_544__96_), .Q(rx_96_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_213 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf1), .D(_544__97_), .Q(rx_97_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_214 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf1), .D(_544__98_), .Q(rx_98_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_215 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf1), .D(_544__99_), .Q(rx_99_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_216 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf1), .D(_544__100_), .Q(rx_100_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_217 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf1), .D(_544__101_), .Q(rx_101_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_218 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf1), .D(_544__102_), .Q(rx_102_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_219 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf1), .D(_544__103_), .Q(rx_103_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_220 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf1), .D(_544__104_), .Q(rx_104_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_221 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf1), .D(_544__105_), .Q(rx_105_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_222 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf1), .D(_544__106_), .Q(rx_106_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_223 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf1), .D(_544__107_), .Q(rx_107_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_224 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__108_), .Q(rx_108_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_225 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__109_), .Q(rx_109_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_226 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf0), .D(_544__110_), .Q(rx_110_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_227 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf0), .D(_544__111_), .Q(rx_111_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_228 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf0), .D(_544__112_), .Q(rx_112_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_229 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf0), .D(_544__113_), .Q(rx_113_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_230 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf0), .D(_544__114_), .Q(rx_114_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_231 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf0), .D(_544__115_), .Q(rx_115_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_232 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf0), .D(_544__116_), .Q(rx_116_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_233 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf0), .D(_544__117_), .Q(rx_117_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_234 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf0), .D(_544__118_), .Q(rx_118_), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_235 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf0), .D(_544__119_), .Q(rx_119_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_236 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf0), .D(_544__120_), .Q(rx_120_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_237 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf0), .D(_544__121_), .Q(rx_121_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_238 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf0), .D(_544__122_), .Q(rx_122_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_239 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf1), .D(_544__123_), .Q(rx_123_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_240 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf0), .D(_544__124_), .Q(rx_124_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_241 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf14_bF_buf3), .D(_544__125_), .Q(rx_125_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_242 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf13_bF_buf3), .D(_544__126_), .Q(rx_126_), .R(_547__bF_buf5), .S(vdd) );
DFFSR DFFSR_243 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf12_bF_buf3), .D(_544__127_), .Q(rx_127_), .R(_547__bF_buf4), .S(vdd) );
DFFSR DFFSR_244 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf11_bF_buf3), .D(_545_), .Q(_423_), .R(_547__bF_buf3), .S(vdd) );
DFFSR DFFSR_245 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf10_bF_buf3), .D(_546_), .Q(clgen_enable), .R(_547__bF_buf2), .S(vdd) );
DFFSR DFFSR_246 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf9_bF_buf3), .D(_543__0_), .Q(shift_cnt_0_), .R(_547__bF_buf1), .S(vdd) );
DFFSR DFFSR_247 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf8_bF_buf3), .D(_543__1_), .Q(shift_cnt_1_), .R(_547__bF_buf0), .S(vdd) );
DFFSR DFFSR_248 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf7_bF_buf3), .D(_543__2_), .Q(shift_cnt_2_), .R(_547__bF_buf10), .S(vdd) );
DFFSR DFFSR_249 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf6_bF_buf3), .D(_543__3_), .Q(shift_cnt_3_), .R(_547__bF_buf9), .S(vdd) );
DFFSR DFFSR_250 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf5_bF_buf3), .D(_543__4_), .Q(shift_cnt_4_), .R(_547__bF_buf8), .S(vdd) );
DFFSR DFFSR_251 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf4_bF_buf3), .D(_543__5_), .Q(shift_cnt_5_), .R(_547__bF_buf7), .S(vdd) );
DFFSR DFFSR_252 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf3_bF_buf3), .D(_543__6_), .Q(shift_cnt_6_), .R(_547__bF_buf6), .S(vdd) );
DFFSR DFFSR_253 ( .gnd(gnd), .vdd(vdd), .CLK(wb_clk_i_bF_buf2_bF_buf3), .D(_543__7_), .Q(shift_cnt_7_), .R(_547__bF_buf5), .S(vdd) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(char_len_0_), .Y(ctrl_0_) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(char_len_1_), .Y(ctrl_1_) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(char_len_2_), .Y(ctrl_2_) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(char_len_3_), .Y(ctrl_3_) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(char_len_4_), .Y(ctrl_4_) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(char_len_5_), .Y(ctrl_5_) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(char_len_6_), .Y(ctrl_6_) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(clgen_go), .Y(ctrl_8_) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(rx_negedge), .Y(ctrl_9_) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(shift_tx_negedge), .Y(ctrl_10_) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(lsb_bF_buf1), .Y(ctrl_11_) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(ie), .Y(ctrl_12_) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(ass), .Y(ctrl_13_) );
endmodule
